VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

SITE CORE_TypTyp_0p4_25
  SYMMETRY y ;
  CLASS core ;
SIZE 0.042 BY 0.384 ; 
END CORE_TypTyp_0p4_25



MACRO AND2_X1
  CLASS core ;
  FOREIGN AND2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.128 0.135 0.348   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.063 0.051 0.262   ; 
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.201 0.057 0.219 0.320   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.177 0.398   ; 
RECT 0.177 0.370 0.259 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.259 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.075 0.081 0.093 0.095   ; 
RECT 0.075 0.095 0.093 0.214   ; 
RECT 0.075 0.214 0.093 0.272   ; 
RECT 0.093 0.081 0.159 0.095   ; 
RECT 0.159 0.081 0.177 0.095   ; 
RECT 0.159 0.095 0.177 0.214   ; 
      LAYER M1 ;
RECT 0.075 0.081 0.093 0.095   ; 
RECT 0.075 0.095 0.093 0.214   ; 
RECT 0.075 0.214 0.093 0.272   ; 
RECT 0.093 0.081 0.159 0.095   ; 
RECT 0.159 0.081 0.177 0.095   ; 
RECT 0.159 0.095 0.177 0.214   ; 
  END
END AND2_X1

MACRO AND2_X2
  CLASS core ;
  FOREIGN AND2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.100 0.128 0.116 0.256   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.025 0.124 0.047 0.260   ; 
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.170 0.032 0.172 0.065   ; 
RECT 0.170 0.319 0.172 0.352   ; 
RECT 0.172 0.032 0.188 0.065   ; 
RECT 0.172 0.065 0.188 0.319   ; 
RECT 0.172 0.319 0.188 0.352   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.006 0.370 0.152 0.398   ; 
RECT 0.152 0.370 0.258 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.006 -0.014 0.258 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.030 0.287 0.046 0.301   ; 
RECT 0.046 0.083 0.136 0.097   ; 
RECT 0.046 0.287 0.136 0.301   ; 
RECT 0.136 0.083 0.152 0.097   ; 
RECT 0.136 0.097 0.152 0.287   ; 
RECT 0.136 0.287 0.152 0.301   ; 
      LAYER M1 ;
RECT 0.030 0.287 0.046 0.301   ; 
RECT 0.046 0.083 0.136 0.097   ; 
RECT 0.046 0.287 0.136 0.301   ; 
RECT 0.136 0.083 0.152 0.097   ; 
RECT 0.136 0.097 0.152 0.287   ; 
RECT 0.136 0.287 0.152 0.301   ; 
  END
END AND2_X2


MACRO AND3_X1
  CLASS core ;
  FOREIGN AND3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.336 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.201 0.096 0.219 0.288   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.113 0.096 0.138 0.288   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.032 0.096 0.052 0.288   ; 
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.285 0.057 0.303 0.327   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.261 0.398   ; 
RECT 0.261 0.370 0.343 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.343 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.052 0.050 0.156 0.066   ; 
RECT 0.035 0.316 0.180 0.330   ; 
RECT 0.180 0.048 0.243 0.068   ; 
RECT 0.180 0.316 0.243 0.330   ; 
RECT 0.243 0.048 0.261 0.068   ; 
RECT 0.243 0.068 0.261 0.316   ; 
RECT 0.243 0.316 0.261 0.330   ; 
      LAYER M1 ;
RECT 0.052 0.050 0.156 0.066   ; 
RECT 0.035 0.316 0.180 0.330   ; 
RECT 0.180 0.048 0.243 0.068   ; 
RECT 0.180 0.316 0.243 0.330   ; 
RECT 0.243 0.048 0.261 0.068   ; 
RECT 0.243 0.068 0.261 0.316   ; 
RECT 0.243 0.316 0.261 0.330   ; 
  END
END AND3_X1

MACRO AND3_X2
  CLASS core ;
  FOREIGN AND3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.336 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.160 0.135 0.256   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.030 0.128 0.054 0.256   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.159 0.151 0.177 0.268   ; 
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.240 0.032 0.243 0.078   ; 
RECT 0.240 0.319 0.243 0.352   ; 
RECT 0.243 0.032 0.261 0.078   ; 
RECT 0.243 0.078 0.261 0.319   ; 
RECT 0.243 0.319 0.261 0.352   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.219 0.398   ; 
RECT 0.219 0.370 0.343 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.343 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.032 0.036 0.052 0.078   ; 
RECT 0.032 0.078 0.052 0.094   ; 
RECT 0.052 0.078 0.196 0.094   ; 
RECT 0.035 0.290 0.096 0.306   ; 
RECT 0.096 0.112 0.201 0.126   ; 
RECT 0.096 0.290 0.201 0.306   ; 
RECT 0.201 0.112 0.219 0.126   ; 
RECT 0.201 0.126 0.219 0.290   ; 
RECT 0.201 0.290 0.219 0.306   ; 
      LAYER M1 ;
RECT 0.032 0.036 0.052 0.078   ; 
RECT 0.032 0.078 0.052 0.094   ; 
RECT 0.052 0.078 0.196 0.094   ; 
RECT 0.035 0.290 0.096 0.306   ; 
RECT 0.096 0.112 0.201 0.126   ; 
RECT 0.096 0.290 0.201 0.306   ; 
RECT 0.201 0.112 0.219 0.126   ; 
RECT 0.201 0.126 0.219 0.290   ; 
RECT 0.201 0.290 0.219 0.306   ; 
  END
END AND3_X2

MACRO AND4_X1
  CLASS core ;
  FOREIGN AND4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.378 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.243 0.096 0.261 0.288   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.158 0.096 0.178 0.288   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.096 0.093 0.256   ; 
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.096 0.051 0.288   ; 
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.327 0.057 0.345 0.327   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.303 0.398   ; 
RECT 0.303 0.370 0.385 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.385 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.054 0.318 0.222 0.334   ; 
RECT 0.222 0.050 0.285 0.066   ; 
RECT 0.222 0.318 0.285 0.334   ; 
RECT 0.285 0.050 0.303 0.066   ; 
RECT 0.285 0.066 0.303 0.318   ; 
RECT 0.285 0.318 0.303 0.334   ; 
RECT 0.092 0.050 0.196 0.074   ; 
      LAYER M1 ;
RECT 0.054 0.318 0.222 0.334   ; 
RECT 0.222 0.050 0.285 0.066   ; 
RECT 0.222 0.318 0.285 0.334   ; 
RECT 0.285 0.050 0.303 0.066   ; 
RECT 0.285 0.066 0.303 0.318   ; 
RECT 0.285 0.318 0.303 0.334   ; 
RECT 0.092 0.050 0.196 0.074   ; 
  END
END AND4_X1

MACRO AND4_X2
  CLASS core ;
  FOREIGN AND4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.378 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.219 0.120 0.235 0.288   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.143 0.096 0.159 0.289   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.067 0.096 0.084 0.289   ; 
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.030 0.096 0.046 0.289   ; 
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.294 0.048 0.311 0.320   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.006 0.370 0.273 0.398   ; 
RECT 0.273 0.370 0.384 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.006 -0.014 0.384 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.084 0.050 0.176 0.066   ; 
RECT 0.048 0.318 0.202 0.334   ; 
RECT 0.202 0.082 0.256 0.098   ; 
RECT 0.202 0.318 0.256 0.334   ; 
RECT 0.256 0.082 0.273 0.098   ; 
RECT 0.256 0.098 0.273 0.318   ; 
RECT 0.256 0.318 0.273 0.334   ; 
      LAYER M1 ;
RECT 0.084 0.050 0.176 0.066   ; 
RECT 0.048 0.318 0.202 0.334   ; 
RECT 0.202 0.082 0.256 0.098   ; 
RECT 0.202 0.318 0.256 0.334   ; 
RECT 0.256 0.082 0.273 0.098   ; 
RECT 0.256 0.098 0.273 0.318   ; 
RECT 0.256 0.318 0.273 0.334   ; 
  END
END AND4_X2

MACRO ANTENNA
  CLASS core ;
  FOREIGN ANTENNA 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.126 BY 0.384 ; 
END ANTENNA

MACRO AOI21_X1
  CLASS core ;
  FOREIGN AOI21_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.096 0.135 0.256   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.067 0.051 0.256   ; 
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.201 0.096 0.219 0.256   ; 
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.050 0.093 0.066   ; 
RECT 0.075 0.066 0.093 0.268   ; 
RECT 0.093 0.050 0.201 0.066   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.196 0.398   ; 
RECT 0.196 0.370 0.259 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.259 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.032 0.290 0.052 0.306   ; 
RECT 0.032 0.306 0.052 0.352   ; 
RECT 0.052 0.290 0.196 0.306   ; 
      LAYER M1 ;
RECT 0.032 0.290 0.052 0.306   ; 
RECT 0.032 0.306 0.052 0.352   ; 
RECT 0.052 0.290 0.196 0.306   ; 
  END
END AOI21_X1

MACRO AOI21_X2
  CLASS core ;
  FOREIGN AOI21_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.162 0.151 0.174 0.224   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.106 0.115 0.118 0.129   ; 
RECT 0.106 0.129 0.118 0.224   ; 
RECT 0.106 0.224 0.118 0.256   ; 
RECT 0.118 0.115 0.216 0.129   ; 
RECT 0.216 0.115 0.232 0.129   ; 
RECT 0.216 0.129 0.232 0.224   ; 
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.050 0.128 0.062 0.224   ; 
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.034 0.083 0.078 0.097   ; 
RECT 0.078 0.083 0.090 0.097   ; 
RECT 0.078 0.097 0.090 0.245   ; 
RECT 0.078 0.245 0.090 0.286   ; 
RECT 0.078 0.286 0.090 0.299   ; 
RECT 0.090 0.083 0.188 0.097   ; 
RECT 0.090 0.286 0.188 0.299   ; 
RECT 0.188 0.286 0.190 0.299   ; 
RECT 0.190 0.245 0.202 0.286   ; 
RECT 0.190 0.286 0.202 0.299   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.370 0.230 0.398   ; 
RECT 0.230 0.370 0.234 0.398   ; 
RECT 0.234 0.370 0.256 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.014 0.256 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.021 0.275 0.035 0.318   ; 
RECT 0.021 0.318 0.035 0.334   ; 
RECT 0.035 0.318 0.218 0.334   ; 
RECT 0.218 0.258 0.230 0.275   ; 
RECT 0.218 0.275 0.230 0.318   ; 
RECT 0.218 0.318 0.230 0.334   ; 
RECT 0.064 0.051 0.234 0.065   ; 
      LAYER M1 ;
RECT 0.021 0.275 0.035 0.318   ; 
RECT 0.021 0.318 0.035 0.334   ; 
RECT 0.035 0.318 0.218 0.334   ; 
RECT 0.218 0.258 0.230 0.275   ; 
RECT 0.218 0.275 0.230 0.318   ; 
RECT 0.218 0.318 0.230 0.334   ; 
RECT 0.064 0.051 0.234 0.065   ; 
  END
END AOI21_X2

MACRO AOI22_X1
  CLASS core ;
  FOREIGN AOI22_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.159 0.096 0.177 0.256   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.243 0.096 0.261 0.242   ; 
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.099 0.093 0.288   ; 
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.096 0.051 0.288   ; 
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.092 0.051 0.201 0.065   ; 
RECT 0.201 0.051 0.219 0.065   ; 
RECT 0.201 0.065 0.219 0.291   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.261 0.398   ; 
RECT 0.261 0.370 0.301 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.301 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.054 0.315 0.243 0.337   ; 
RECT 0.243 0.276 0.261 0.315   ; 
RECT 0.243 0.315 0.261 0.337   ; 
      LAYER M1 ;
RECT 0.054 0.315 0.243 0.337   ; 
RECT 0.243 0.276 0.261 0.315   ; 
RECT 0.243 0.315 0.261 0.337   ; 
  END
END AOI22_X1

MACRO AOI22_X2
  CLASS core ;
  FOREIGN AOI22_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.166 0.137 0.177 0.151   ; 
RECT 0.166 0.151 0.177 0.245   ; 
RECT 0.166 0.245 0.177 0.256   ; 
RECT 0.177 0.137 0.250 0.151   ; 
RECT 0.250 0.137 0.264 0.151   ; 
RECT 0.264 0.137 0.275 0.151   ; 
RECT 0.264 0.151 0.275 0.245   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.215 0.185 0.226 0.256   ; 
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.153 0.128 0.263   ; 
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.019 0.121 0.030 0.256   ; 
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.093 0.100 0.103 0.114   ; 
RECT 0.093 0.114 0.103 0.114   ; 
RECT 0.093 0.114 0.103 0.160   ; 
RECT 0.103 0.100 0.139 0.114   ; 
RECT 0.139 0.100 0.142 0.114   ; 
RECT 0.142 0.100 0.152 0.114   ; 
RECT 0.142 0.114 0.152 0.114   ; 
RECT 0.142 0.114 0.152 0.160   ; 
RECT 0.142 0.160 0.152 0.232   ; 
RECT 0.142 0.232 0.152 0.284   ; 
RECT 0.142 0.284 0.152 0.301   ; 
RECT 0.152 0.100 0.240 0.114   ; 
RECT 0.152 0.114 0.240 0.114   ; 
RECT 0.152 0.284 0.240 0.301   ; 
RECT 0.240 0.100 0.250 0.114   ; 
RECT 0.240 0.114 0.250 0.114   ; 
RECT 0.240 0.232 0.250 0.284   ; 
RECT 0.240 0.284 0.250 0.301   ; 
RECT 0.250 0.100 0.264 0.114   ; 
RECT 0.250 0.114 0.264 0.114   ; 
RECT 0.264 0.048 0.275 0.100   ; 
RECT 0.264 0.100 0.275 0.114   ; 
RECT 0.264 0.114 0.275 0.114   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.370 0.275 0.398   ; 
RECT 0.275 0.370 0.298 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.014 0.298 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.155 0.066 0.240 0.082   ; 
RECT 0.240 0.036 0.250 0.066   ; 
RECT 0.240 0.066 0.250 0.082   ; 
RECT 0.029 0.319 0.264 0.333   ; 
RECT 0.264 0.279 0.275 0.319   ; 
RECT 0.264 0.319 0.275 0.333   ; 
RECT 0.033 0.043 0.139 0.072   ; 
      LAYER M1 ;
RECT 0.155 0.066 0.240 0.082   ; 
RECT 0.240 0.036 0.250 0.066   ; 
RECT 0.240 0.066 0.250 0.082   ; 
RECT 0.029 0.319 0.264 0.333   ; 
RECT 0.264 0.279 0.275 0.319   ; 
RECT 0.264 0.319 0.275 0.333   ; 
RECT 0.033 0.043 0.139 0.072   ; 
  END
END AOI22_X2

MACRO BUF_X1
  CLASS core ;
  FOREIGN BUF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.210 BY 0.384 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.096 0.051 0.288   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.158 0.057 0.178 0.352   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.094 0.398   ; 
RECT 0.094 0.370 0.217 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.217 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.075 0.036 0.075 0.092   ; 
RECT 0.075 0.092 0.075 0.106   ; 
RECT 0.075 0.214 0.075 0.228   ; 
RECT 0.075 0.228 0.075 0.279   ; 
RECT 0.075 0.036 0.093 0.092   ; 
RECT 0.075 0.092 0.093 0.106   ; 
RECT 0.075 0.106 0.093 0.214   ; 
RECT 0.075 0.214 0.093 0.228   ; 
RECT 0.075 0.228 0.093 0.279   ; 
RECT 0.093 0.092 0.094 0.106   ; 
RECT 0.093 0.106 0.094 0.214   ; 
RECT 0.093 0.214 0.094 0.228   ; 
      LAYER M1 ;
RECT 0.075 0.036 0.075 0.092   ; 
RECT 0.075 0.092 0.075 0.106   ; 
RECT 0.075 0.214 0.075 0.228   ; 
RECT 0.075 0.228 0.075 0.279   ; 
RECT 0.075 0.036 0.093 0.092   ; 
RECT 0.075 0.092 0.093 0.106   ; 
RECT 0.075 0.106 0.093 0.214   ; 
RECT 0.075 0.214 0.093 0.228   ; 
RECT 0.075 0.228 0.093 0.279   ; 
RECT 0.093 0.092 0.094 0.106   ; 
RECT 0.093 0.106 0.094 0.214   ; 
RECT 0.093 0.214 0.094 0.228   ; 
  END
END BUF_X1

MACRO BUF_X2
  CLASS core ;
  FOREIGN BUF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.210 BY 0.384 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.134 0.051 0.256   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.114 0.302 0.116 0.352   ; 
RECT 0.116 0.036 0.117 0.066   ; 
RECT 0.116 0.302 0.117 0.352   ; 
RECT 0.117 0.036 0.135 0.066   ; 
RECT 0.117 0.066 0.135 0.302   ; 
RECT 0.117 0.302 0.135 0.352   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.093 0.398   ; 
RECT 0.093 0.370 0.217 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.217 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.028 0.278 0.033 0.292   ; 
RECT 0.028 0.292 0.033 0.343   ; 
RECT 0.033 0.048 0.051 0.096   ; 
RECT 0.033 0.096 0.051 0.110   ; 
RECT 0.033 0.278 0.051 0.292   ; 
RECT 0.033 0.292 0.051 0.343   ; 
RECT 0.051 0.096 0.056 0.110   ; 
RECT 0.051 0.278 0.056 0.292   ; 
RECT 0.051 0.292 0.056 0.343   ; 
RECT 0.056 0.096 0.075 0.110   ; 
RECT 0.056 0.278 0.075 0.292   ; 
RECT 0.075 0.096 0.093 0.110   ; 
RECT 0.075 0.110 0.093 0.278   ; 
RECT 0.075 0.278 0.093 0.292   ; 
      LAYER M1 ;
RECT 0.028 0.278 0.033 0.292   ; 
RECT 0.028 0.292 0.033 0.343   ; 
RECT 0.033 0.048 0.051 0.096   ; 
RECT 0.033 0.096 0.051 0.110   ; 
RECT 0.033 0.278 0.051 0.292   ; 
RECT 0.033 0.292 0.051 0.343   ; 
RECT 0.051 0.096 0.056 0.110   ; 
RECT 0.051 0.278 0.056 0.292   ; 
RECT 0.051 0.292 0.056 0.343   ; 
RECT 0.056 0.096 0.075 0.110   ; 
RECT 0.056 0.278 0.075 0.292   ; 
RECT 0.075 0.096 0.093 0.110   ; 
RECT 0.075 0.110 0.093 0.278   ; 
RECT 0.075 0.278 0.093 0.292   ; 
  END
END BUF_X2

MACRO BUF_X4
  CLASS core ;
  FOREIGN BUF_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.210 BY 0.384 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.073 0.121 0.084 0.263   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.059 0.051 0.086 0.065   ; 
RECT 0.086 0.051 0.111 0.065   ; 
RECT 0.086 0.319 0.111 0.333   ; 
RECT 0.111 0.051 0.151 0.065   ; 
RECT 0.111 0.319 0.151 0.333   ; 
RECT 0.151 0.051 0.164 0.065   ; 
RECT 0.151 0.065 0.164 0.319   ; 
RECT 0.151 0.319 0.164 0.333   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.370 0.111 0.398   ; 
RECT 0.111 0.370 0.214 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.014 0.214 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.011 0.083 0.035 0.099   ; 
RECT 0.035 0.083 0.099 0.099   ; 
RECT 0.035 0.285 0.099 0.301   ; 
RECT 0.099 0.083 0.111 0.099   ; 
RECT 0.099 0.099 0.111 0.285   ; 
RECT 0.099 0.285 0.111 0.301   ; 
      LAYER M1 ;
RECT 0.011 0.083 0.035 0.099   ; 
RECT 0.035 0.083 0.099 0.099   ; 
RECT 0.035 0.285 0.099 0.301   ; 
RECT 0.099 0.083 0.111 0.099   ; 
RECT 0.099 0.099 0.111 0.285   ; 
RECT 0.099 0.285 0.111 0.301   ; 
  END
END BUF_X4

MACRO BUF_X8
  CLASS core ;
  FOREIGN BUF_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.210 BY 0.384 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.012 0.128 0.018 0.183   ; 
RECT 0.012 0.183 0.018 0.199   ; 
RECT 0.012 0.199 0.018 0.256   ; 
RECT 0.018 0.183 0.070 0.199   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.079 0.051 0.164 0.065   ; 
RECT 0.079 0.319 0.164 0.333   ; 
RECT 0.164 0.051 0.177 0.065   ; 
RECT 0.164 0.319 0.177 0.333   ; 
RECT 0.177 0.051 0.183 0.065   ; 
RECT 0.177 0.065 0.183 0.319   ; 
RECT 0.177 0.319 0.183 0.333   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 0.370 0.164 0.398   ; 
RECT 0.164 0.370 0.212 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 -0.014 0.212 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.023 0.049 0.027 0.093   ; 
RECT 0.023 0.093 0.027 0.107   ; 
RECT 0.027 0.049 0.033 0.093   ; 
RECT 0.027 0.093 0.033 0.107   ; 
RECT 0.027 0.264 0.033 0.292   ; 
RECT 0.027 0.292 0.033 0.335   ; 
RECT 0.033 0.049 0.037 0.093   ; 
RECT 0.033 0.093 0.037 0.107   ; 
RECT 0.033 0.264 0.037 0.292   ; 
RECT 0.037 0.093 0.083 0.107   ; 
RECT 0.037 0.264 0.083 0.292   ; 
RECT 0.083 0.093 0.090 0.107   ; 
RECT 0.083 0.107 0.090 0.171   ; 
RECT 0.083 0.171 0.090 0.184   ; 
RECT 0.083 0.184 0.090 0.264   ; 
RECT 0.083 0.264 0.090 0.292   ; 
RECT 0.090 0.171 0.164 0.184   ; 
      LAYER M1 ;
RECT 0.023 0.049 0.027 0.093   ; 
RECT 0.023 0.093 0.027 0.107   ; 
RECT 0.027 0.049 0.033 0.093   ; 
RECT 0.027 0.093 0.033 0.107   ; 
RECT 0.027 0.264 0.033 0.292   ; 
RECT 0.027 0.292 0.033 0.335   ; 
RECT 0.033 0.049 0.037 0.093   ; 
RECT 0.033 0.093 0.037 0.107   ; 
RECT 0.033 0.264 0.037 0.292   ; 
RECT 0.037 0.093 0.083 0.107   ; 
RECT 0.037 0.264 0.083 0.292   ; 
RECT 0.083 0.093 0.090 0.107   ; 
RECT 0.083 0.107 0.090 0.171   ; 
RECT 0.083 0.171 0.090 0.184   ; 
RECT 0.083 0.184 0.090 0.264   ; 
RECT 0.083 0.264 0.090 0.292   ; 
RECT 0.090 0.171 0.164 0.184   ; 
  END
END BUF_X8

MACRO BUF_X12
  CLASS core ;
  FOREIGN BUF_X12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.384 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.010 0.118 0.017 0.183   ; 
RECT 0.010 0.183 0.017 0.199   ; 
RECT 0.010 0.199 0.017 0.258   ; 
RECT 0.017 0.183 0.093 0.199   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.102 0.051 0.234 0.065   ; 
RECT 0.102 0.319 0.234 0.333   ; 
RECT 0.234 0.051 0.248 0.065   ; 
RECT 0.234 0.319 0.248 0.333   ; 
RECT 0.248 0.051 0.255 0.065   ; 
RECT 0.248 0.065 0.255 0.319   ; 
RECT 0.248 0.319 0.255 0.333   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 0.370 0.234 0.398   ; 
RECT 0.234 0.370 0.282 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 -0.014 0.282 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.021 0.276 0.024 0.292   ; 
RECT 0.021 0.292 0.024 0.335   ; 
RECT 0.024 0.049 0.031 0.092   ; 
RECT 0.024 0.092 0.031 0.108   ; 
RECT 0.024 0.276 0.031 0.292   ; 
RECT 0.024 0.292 0.031 0.335   ; 
RECT 0.031 0.092 0.034 0.108   ; 
RECT 0.031 0.276 0.034 0.292   ; 
RECT 0.031 0.292 0.034 0.335   ; 
RECT 0.034 0.092 0.101 0.108   ; 
RECT 0.034 0.276 0.101 0.292   ; 
RECT 0.101 0.092 0.107 0.108   ; 
RECT 0.101 0.108 0.107 0.185   ; 
RECT 0.101 0.185 0.107 0.199   ; 
RECT 0.101 0.199 0.107 0.276   ; 
RECT 0.101 0.276 0.107 0.292   ; 
RECT 0.107 0.185 0.234 0.199   ; 
      LAYER M1 ;
RECT 0.021 0.276 0.024 0.292   ; 
RECT 0.021 0.292 0.024 0.335   ; 
RECT 0.024 0.049 0.031 0.092   ; 
RECT 0.024 0.092 0.031 0.108   ; 
RECT 0.024 0.276 0.031 0.292   ; 
RECT 0.024 0.292 0.031 0.335   ; 
RECT 0.031 0.092 0.034 0.108   ; 
RECT 0.031 0.276 0.034 0.292   ; 
RECT 0.031 0.292 0.034 0.335   ; 
RECT 0.034 0.092 0.101 0.108   ; 
RECT 0.034 0.276 0.101 0.292   ; 
RECT 0.101 0.092 0.107 0.108   ; 
RECT 0.101 0.108 0.107 0.185   ; 
RECT 0.101 0.185 0.107 0.199   ; 
RECT 0.101 0.199 0.107 0.276   ; 
RECT 0.101 0.276 0.107 0.292   ; 
RECT 0.107 0.185 0.234 0.199   ; 
  END
END BUF_X12


MACRO BUF_X16
  CLASS core ;
  FOREIGN BUF_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.384 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.008 0.116 0.013 0.178   ; 
RECT 0.008 0.178 0.013 0.206   ; 
RECT 0.008 0.206 0.013 0.256   ; 
RECT 0.013 0.178 0.093 0.206   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.100 0.051 0.245 0.065   ; 
RECT 0.100 0.316 0.245 0.330   ; 
RECT 0.245 0.051 0.256 0.065   ; 
RECT 0.245 0.316 0.256 0.330   ; 
RECT 0.256 0.051 0.261 0.065   ; 
RECT 0.256 0.065 0.261 0.316   ; 
RECT 0.256 0.316 0.261 0.330   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 0.370 0.245 0.398   ; 
RECT 0.245 0.370 0.282 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 -0.014 0.282 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.019 0.049 0.024 0.103   ; 
RECT 0.019 0.103 0.024 0.117   ; 
RECT 0.019 0.229 0.024 0.243   ; 
RECT 0.019 0.243 0.024 0.322   ; 
RECT 0.024 0.103 0.099 0.117   ; 
RECT 0.024 0.229 0.099 0.243   ; 
RECT 0.099 0.103 0.104 0.117   ; 
RECT 0.099 0.117 0.104 0.184   ; 
RECT 0.099 0.184 0.104 0.198   ; 
RECT 0.099 0.198 0.104 0.229   ; 
RECT 0.099 0.229 0.104 0.243   ; 
RECT 0.104 0.184 0.245 0.198   ; 
      LAYER M1 ;
RECT 0.019 0.049 0.024 0.103   ; 
RECT 0.019 0.103 0.024 0.117   ; 
RECT 0.019 0.229 0.024 0.243   ; 
RECT 0.019 0.243 0.024 0.322   ; 
RECT 0.024 0.103 0.099 0.117   ; 
RECT 0.024 0.229 0.099 0.243   ; 
RECT 0.099 0.103 0.104 0.117   ; 
RECT 0.099 0.117 0.104 0.184   ; 
RECT 0.099 0.184 0.104 0.198   ; 
RECT 0.099 0.198 0.104 0.229   ; 
RECT 0.099 0.229 0.104 0.243   ; 
RECT 0.104 0.184 0.245 0.198   ; 
  END
END BUF_X16

MACRO CLKBUF_X1
  CLASS core ;
  FOREIGN CLKBUF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.210 BY 0.384 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.096 0.051 0.288   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.158 0.057 0.178 0.352   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.094 0.398   ; 
RECT 0.094 0.370 0.217 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.217 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.075 0.036 0.075 0.092   ; 
RECT 0.075 0.092 0.075 0.106   ; 
RECT 0.075 0.196 0.075 0.229   ; 
RECT 0.075 0.229 0.075 0.262   ; 
RECT 0.075 0.036 0.093 0.092   ; 
RECT 0.075 0.092 0.093 0.106   ; 
RECT 0.075 0.106 0.093 0.196   ; 
RECT 0.075 0.196 0.093 0.229   ; 
RECT 0.075 0.229 0.093 0.262   ; 
RECT 0.093 0.092 0.094 0.106   ; 
RECT 0.093 0.106 0.094 0.196   ; 
RECT 0.093 0.196 0.094 0.229   ; 
      LAYER M1 ;
RECT 0.075 0.036 0.075 0.092   ; 
RECT 0.075 0.092 0.075 0.106   ; 
RECT 0.075 0.196 0.075 0.229   ; 
RECT 0.075 0.229 0.075 0.262   ; 
RECT 0.075 0.036 0.093 0.092   ; 
RECT 0.075 0.092 0.093 0.106   ; 
RECT 0.075 0.106 0.093 0.196   ; 
RECT 0.075 0.196 0.093 0.229   ; 
RECT 0.075 0.229 0.093 0.262   ; 
RECT 0.093 0.092 0.094 0.106   ; 
RECT 0.093 0.106 0.094 0.196   ; 
RECT 0.093 0.196 0.094 0.229   ; 
  END
END CLKBUF_X1

MACRO CLKBUF_X2
  CLASS core ;
  FOREIGN CLKBUF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.210 BY 0.384 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.148 0.051 0.256   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.114 0.319 0.117 0.352   ; 
RECT 0.117 0.036 0.135 0.319   ; 
RECT 0.117 0.319 0.135 0.352   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.093 0.398   ; 
RECT 0.093 0.370 0.217 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.217 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.032 0.065 0.052 0.096   ; 
RECT 0.032 0.096 0.052 0.110   ; 
RECT 0.032 0.278 0.052 0.292   ; 
RECT 0.032 0.292 0.052 0.343   ; 
RECT 0.052 0.096 0.075 0.110   ; 
RECT 0.052 0.278 0.075 0.292   ; 
RECT 0.075 0.096 0.093 0.110   ; 
RECT 0.075 0.110 0.093 0.278   ; 
RECT 0.075 0.278 0.093 0.292   ; 
      LAYER M1 ;
RECT 0.032 0.065 0.052 0.096   ; 
RECT 0.032 0.096 0.052 0.110   ; 
RECT 0.032 0.278 0.052 0.292   ; 
RECT 0.032 0.292 0.052 0.343   ; 
RECT 0.052 0.096 0.075 0.110   ; 
RECT 0.052 0.278 0.075 0.292   ; 
RECT 0.075 0.096 0.093 0.110   ; 
RECT 0.075 0.110 0.093 0.278   ; 
RECT 0.075 0.278 0.093 0.292   ; 
  END
END CLKBUF_X2

MACRO CLKBUF_X4
  CLASS core ;
  FOREIGN CLKBUF_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.210 BY 0.384 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.047 0.121 0.058 0.263   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.059 0.051 0.084 0.065   ; 
RECT 0.084 0.051 0.084 0.065   ; 
RECT 0.084 0.319 0.084 0.333   ; 
RECT 0.084 0.051 0.151 0.065   ; 
RECT 0.084 0.319 0.151 0.333   ; 
RECT 0.151 0.051 0.164 0.065   ; 
RECT 0.151 0.065 0.164 0.319   ; 
RECT 0.151 0.319 0.164 0.333   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.370 0.084 0.398   ; 
RECT 0.084 0.370 0.214 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.014 0.214 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.017 0.083 0.034 0.097   ; 
RECT 0.034 0.083 0.073 0.097   ; 
RECT 0.034 0.287 0.073 0.301   ; 
RECT 0.073 0.083 0.084 0.097   ; 
RECT 0.073 0.097 0.084 0.287   ; 
RECT 0.073 0.287 0.084 0.301   ; 
      LAYER M1 ;
RECT 0.017 0.083 0.034 0.097   ; 
RECT 0.034 0.083 0.073 0.097   ; 
RECT 0.034 0.287 0.073 0.301   ; 
RECT 0.073 0.083 0.084 0.097   ; 
RECT 0.073 0.097 0.084 0.287   ; 
RECT 0.073 0.287 0.084 0.301   ; 
  END
END CLKBUF_X4

MACRO CLKBUF_X8
  CLASS core ;
  FOREIGN CLKBUF_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.210 BY 0.384 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.012 0.128 0.018 0.164   ; 
RECT 0.012 0.164 0.018 0.178   ; 
RECT 0.012 0.178 0.018 0.256   ; 
RECT 0.018 0.128 0.019 0.164   ; 
RECT 0.018 0.164 0.019 0.178   ; 
RECT 0.019 0.164 0.075 0.178   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.079 0.051 0.168 0.065   ; 
RECT 0.079 0.319 0.168 0.333   ; 
RECT 0.168 0.051 0.177 0.065   ; 
RECT 0.168 0.319 0.177 0.333   ; 
RECT 0.177 0.051 0.183 0.065   ; 
RECT 0.177 0.065 0.183 0.319   ; 
RECT 0.177 0.319 0.183 0.333   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 0.370 0.168 0.398   ; 
RECT 0.168 0.370 0.212 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 -0.014 0.212 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.012 0.083 0.027 0.097   ; 
RECT 0.027 0.083 0.033 0.097   ; 
RECT 0.027 0.225 0.033 0.241   ; 
RECT 0.027 0.241 0.033 0.271   ; 
RECT 0.033 0.083 0.095 0.097   ; 
RECT 0.033 0.225 0.095 0.241   ; 
RECT 0.095 0.083 0.102 0.097   ; 
RECT 0.095 0.097 0.102 0.178   ; 
RECT 0.095 0.178 0.102 0.207   ; 
RECT 0.095 0.207 0.102 0.225   ; 
RECT 0.095 0.225 0.102 0.241   ; 
RECT 0.102 0.178 0.168 0.207   ; 
      LAYER M1 ;
RECT 0.012 0.083 0.027 0.097   ; 
RECT 0.027 0.083 0.033 0.097   ; 
RECT 0.027 0.225 0.033 0.241   ; 
RECT 0.027 0.241 0.033 0.271   ; 
RECT 0.033 0.083 0.095 0.097   ; 
RECT 0.033 0.225 0.095 0.241   ; 
RECT 0.095 0.083 0.102 0.097   ; 
RECT 0.095 0.097 0.102 0.178   ; 
RECT 0.095 0.178 0.102 0.207   ; 
RECT 0.095 0.207 0.102 0.225   ; 
RECT 0.095 0.225 0.102 0.241   ; 
RECT 0.102 0.178 0.168 0.207   ; 
  END
END CLKBUF_X8

MACRO CLKBUF_X12
  CLASS core ;
  FOREIGN CLKBUF_X12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.384 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.010 0.119 0.018 0.168   ; 
RECT 0.010 0.168 0.018 0.184   ; 
RECT 0.010 0.184 0.018 0.265   ; 
RECT 0.018 0.168 0.093 0.184   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.102 0.051 0.218 0.065   ; 
RECT 0.102 0.319 0.218 0.333   ; 
RECT 0.218 0.051 0.248 0.065   ; 
RECT 0.218 0.319 0.248 0.333   ; 
RECT 0.248 0.051 0.255 0.065   ; 
RECT 0.248 0.065 0.255 0.319   ; 
RECT 0.248 0.319 0.255 0.333   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 0.370 0.218 0.398   ; 
RECT 0.218 0.370 0.282 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 -0.014 0.282 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.009 0.083 0.025 0.097   ; 
RECT 0.025 0.083 0.031 0.097   ; 
RECT 0.025 0.275 0.031 0.289   ; 
RECT 0.025 0.289 0.031 0.335   ; 
RECT 0.031 0.083 0.101 0.097   ; 
RECT 0.031 0.275 0.101 0.289   ; 
RECT 0.101 0.083 0.107 0.097   ; 
RECT 0.101 0.097 0.107 0.157   ; 
RECT 0.101 0.157 0.107 0.173   ; 
RECT 0.101 0.173 0.107 0.275   ; 
RECT 0.101 0.275 0.107 0.289   ; 
RECT 0.107 0.083 0.108 0.097   ; 
RECT 0.107 0.097 0.108 0.157   ; 
RECT 0.107 0.157 0.108 0.173   ; 
RECT 0.108 0.157 0.218 0.173   ; 
      LAYER M1 ;
RECT 0.009 0.083 0.025 0.097   ; 
RECT 0.025 0.083 0.031 0.097   ; 
RECT 0.025 0.275 0.031 0.289   ; 
RECT 0.025 0.289 0.031 0.335   ; 
RECT 0.031 0.083 0.101 0.097   ; 
RECT 0.031 0.275 0.101 0.289   ; 
RECT 0.101 0.083 0.107 0.097   ; 
RECT 0.101 0.097 0.107 0.157   ; 
RECT 0.101 0.157 0.107 0.173   ; 
RECT 0.101 0.173 0.107 0.275   ; 
RECT 0.101 0.275 0.107 0.289   ; 
RECT 0.107 0.083 0.108 0.097   ; 
RECT 0.107 0.097 0.108 0.157   ; 
RECT 0.107 0.157 0.108 0.173   ; 
RECT 0.108 0.157 0.218 0.173   ; 
  END
END CLKBUF_X12

MACRO CLKBUF_X16
  CLASS core ;
  FOREIGN CLKBUF_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.384 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.008 0.111 0.013 0.163   ; 
RECT 0.008 0.163 0.013 0.179   ; 
RECT 0.008 0.179 0.013 0.263   ; 
RECT 0.013 0.163 0.093 0.179   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.100 0.043 0.245 0.072   ; 
RECT 0.100 0.312 0.245 0.341   ; 
RECT 0.245 0.043 0.256 0.072   ; 
RECT 0.245 0.312 0.256 0.341   ; 
RECT 0.256 0.043 0.261 0.072   ; 
RECT 0.256 0.072 0.261 0.312   ; 
RECT 0.256 0.312 0.261 0.341   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 0.370 0.245 0.398   ; 
RECT 0.245 0.370 0.282 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 -0.014 0.282 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.019 0.055 0.024 0.103   ; 
RECT 0.019 0.103 0.024 0.117   ; 
RECT 0.019 0.263 0.024 0.281   ; 
RECT 0.019 0.281 0.024 0.319   ; 
RECT 0.024 0.103 0.100 0.117   ; 
RECT 0.024 0.263 0.100 0.281   ; 
RECT 0.100 0.103 0.110 0.117   ; 
RECT 0.100 0.117 0.110 0.158   ; 
RECT 0.100 0.158 0.110 0.172   ; 
RECT 0.100 0.172 0.110 0.263   ; 
RECT 0.100 0.263 0.110 0.281   ; 
RECT 0.110 0.158 0.245 0.172   ; 
      LAYER M1 ;
RECT 0.019 0.055 0.024 0.103   ; 
RECT 0.019 0.103 0.024 0.117   ; 
RECT 0.019 0.263 0.024 0.281   ; 
RECT 0.019 0.281 0.024 0.319   ; 
RECT 0.024 0.103 0.100 0.117   ; 
RECT 0.024 0.263 0.100 0.281   ; 
RECT 0.100 0.103 0.110 0.117   ; 
RECT 0.100 0.117 0.110 0.158   ; 
RECT 0.100 0.158 0.110 0.172   ; 
RECT 0.100 0.172 0.110 0.263   ; 
RECT 0.100 0.263 0.110 0.281   ; 
RECT 0.110 0.158 0.245 0.172   ; 
  END
END CLKBUF_X16

MACRO DFFRNQ_X1
  CLASS core ;
  FOREIGN DFFRNQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 1.092 BY 0.384 ;

  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 0.149 0.121 0.171 0.263 ;  
    END
  END D

  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
      RECT 0.462 0.156 0.744 0.180 ;  
      RECT 0.744 0.156 0.870 0.180 ;  
    END
  END RN

  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
      RECT 0.021 0.128 0.043 0.256 ;  
    END
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT 1.045 0.032 1.067 0.352 ;  
    END
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT -0.007 0.370 0.093 0.398 ;
      RECT 0.093 0.370 0.135 0.398 ;
      RECT 0.135 0.370 0.219 0.398 ;
      RECT 0.219 0.370 0.261 0.398 ;
      RECT 0.261 0.370 0.345 0.398 ;
      RECT 0.345 0.370 0.534 0.398 ;
      RECT 0.534 0.370 0.597 0.398 ;
      RECT 0.597 0.370 0.639 0.398 ;
      RECT 0.639 0.370 0.723 0.398 ;
      RECT 0.723 0.370 0.780 0.398 ;
      RECT 0.780 0.370 0.977 0.398 ;
      RECT 0.977 0.370 1.099 0.398 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT -0.007 -0.014 1.099 0.014 ;
    END
  END VSS

  OBS
    LAYER MINT1 ;
      RECT 0.0958125 0.137812 0.744125 0.156187 ;
      RECT 0.0538125 0.347813 0.744125 0.366187 ;
    LAYER MINT1 ;
      RECT 0.0958125 0.137812 0.744125 0.156187 ;
      RECT 0.0538125 0.347813 0.744125 0.366187 ;
    LAYER M1 ;
      RECT 0.117 0.036 0.135 0.348 ;
      RECT 0.201 0.036 0.219 0.348 ;
      RECT 0.348 0.312 0.534 0.340 ;
      RECT 0.285 0.051 0.303 0.065 ;
      RECT 0.285 0.065 0.303 0.219 ;
      RECT 0.285 0.219 0.303 0.335 ;
      RECT 0.303 0.051 0.525 0.065 ;
      RECT 0.525 0.051 0.543 0.065 ;
      RECT 0.525 0.065 0.543 0.219 ;
      RECT 0.378 0.165 0.396 0.253 ;
      RECT 0.378 0.253 0.396 0.267 ;
      RECT 0.396 0.253 0.579 0.267 ;
      RECT 0.579 0.036 0.597 0.165 ;
      RECT 0.579 0.165 0.597 0.253 ;
      RECT 0.579 0.253 0.579 0.267 ;
      RECT 0.579 0.267 0.597 0.336 ;
      RECT 0.663 0.051 0.681 0.065 ;
      RECT 0.663 0.065 0.681 0.183 ;
      RECT 0.663 0.183 0.681 0.335 ;
      RECT 0.681 0.051 0.876 0.065 ;
      RECT 0.876 0.051 0.894 0.065 ;
      RECT 0.876 0.065 0.894 0.183 ;
      RECT 0.803 0.197 0.822 0.319 ;
      RECT 0.803 0.319 0.822 0.333 ;
      RECT 0.822 0.319 0.957 0.333 ;
      RECT 0.957 0.036 0.975 0.066 ;
      RECT 0.957 0.066 0.975 0.197 ;
      RECT 0.957 0.197 0.975 0.319 ;
      RECT 0.957 0.319 0.975 0.333 ;
      RECT 0.975 0.066 0.977 0.197 ;
      RECT 0.975 0.197 0.977 0.319 ;
      RECT 0.975 0.319 0.977 0.333 ;
      RECT 0.032 0.042 0.052 0.070 ;
      RECT 0.032 0.070 0.052 0.084 ;
      RECT 0.032 0.283 0.052 0.303 ;
      RECT 0.032 0.303 0.052 0.343 ;
      RECT 0.052 0.070 0.075 0.084 ;
      RECT 0.052 0.283 0.075 0.303 ;
      RECT 0.075 0.070 0.093 0.084 ;
      RECT 0.075 0.084 0.093 0.283 ;
      RECT 0.075 0.283 0.093 0.303 ;
      RECT 0.243 0.097 0.261 0.247 ;
      RECT 0.327 0.201 0.345 0.287 ;
      RECT 0.345 0.097 0.366 0.147 ;
      RECT 0.483 0.129 0.501 0.219 ;
      RECT 0.621 0.137 0.639 0.289 ;
      RECT 0.705 0.087 0.723 0.158 ;
      RECT 0.705 0.230 0.723 0.311 ;
      RECT 0.759 0.083 0.780 0.343 ;
      RECT 0.831 0.087 0.849 0.159 ;
    LAYER V1 ;
      RECT 0.075 0.265 0.093 0.279 ;
      RECT 0.117 0.105 0.135 0.119 ;
      RECT 0.243 0.105 0.261 0.119 ;
      RECT 0.327 0.265 0.345 0.279 ;
      RECT 0.348 0.105 0.366 0.119 ;
      RECT 0.483 0.137 0.501 0.151 ;
      RECT 0.621 0.265 0.639 0.279 ;
      RECT 0.705 0.105 0.723 0.119 ;
      RECT 0.705 0.265 0.723 0.279 ;
      RECT 0.831 0.137 0.849 0.151 ;
    LAYER M1 ;
      RECT 0.117 0.036 0.135 0.348 ;
      RECT 0.201 0.036 0.219 0.348 ;
      RECT 0.348 0.312 0.534 0.340 ;
      RECT 0.285 0.051 0.303 0.065 ;
      RECT 0.285 0.065 0.303 0.219 ;
      RECT 0.285 0.219 0.303 0.335 ;
      RECT 0.303 0.051 0.525 0.065 ;
      RECT 0.525 0.051 0.543 0.065 ;
      RECT 0.525 0.065 0.543 0.219 ;
      RECT 0.378 0.165 0.396 0.253 ;
      RECT 0.378 0.253 0.396 0.267 ;
      RECT 0.396 0.253 0.579 0.267 ;
      RECT 0.579 0.036 0.597 0.165 ;
      RECT 0.579 0.165 0.597 0.253 ;
      RECT 0.579 0.253 0.579 0.267 ;
      RECT 0.579 0.267 0.579 0.336 ;
      RECT 0.663 0.051 0.681 0.065 ;
      RECT 0.663 0.065 0.681 0.183 ;
      RECT 0.663 0.183 0.681 0.335 ;
      RECT 0.681 0.051 0.876 0.065 ;
      RECT 0.876 0.051 0.894 0.065 ;
      RECT 0.876 0.065 0.894 0.183 ;
      RECT 0.803 0.197 0.822 0.319 ;
      RECT 0.803 0.319 0.822 0.333 ;
      RECT 0.822 0.319 0.957 0.333 ;
      RECT 0.957 0.036 0.975 0.066 ;
      RECT 0.957 0.066 0.975 0.197 ;
      RECT 0.957 0.197 0.975 0.319 ;
      RECT 0.957 0.319 0.975 0.333 ;
      RECT 0.975 0.066 0.977 0.197 ;
      RECT 0.975 0.197 0.977 0.319 ;
      RECT 0.975 0.319 0.977 0.333 ;
      RECT 0.032 0.042 0.052 0.070 ;
      RECT 0.032 0.070 0.052 0.084 ;
      RECT 0.032 0.283 0.052 0.303 ;
      RECT 0.032 0.303 0.052 0.343 ;
      RECT 0.052 0.070 0.075 0.084 ;
      RECT 0.052 0.283 0.075 0.303 ;
      RECT 0.075 0.070 0.093 0.084 ;
      RECT 0.075 0.084 0.093 0.283 ;
      RECT 0.075 0.283 0.093 0.303 ;
      RECT 0.243 0.097 0.261 0.247 ;
      RECT 0.327 0.201 0.345 0.287 ;
      RECT 0.345 0.097 0.366 0.147 ;
      RECT 0.483 0.129 0.501 0.219 ;
      RECT 0.621 0.137 0.639 0.289 ;
      RECT 0.705 0.087 0.723 0.158 ;
      RECT 0.705 0.230 0.723 0.311 ;
      RECT 0.759 0.083 0.780 0.343 ;
      RECT 0.831 0.087 0.849 0.159 ;
  END
END DFFRNQ_X1
MACRO DFFSNQ_X1
  CLASS core ;
  FOREIGN DFFSNQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 1.092 BY 0.768 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 0.149 0.159 0.171 0.345 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
      RECT 0.474 0.156 0.744 0.180 ;
      RECT 0.744 0.156 0.870 0.180 ;
    END
  END SN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
      RECT 0.021 0.168 0.043 0.336 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT 1.045 0.042 1.067 0.462 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT -0.007 0.486 0.093 0.522 ;
      RECT 0.093 0.486 0.135 0.522 ;
      RECT 0.135 0.486 0.219 0.522 ;
      RECT 0.219 0.486 0.261 0.522 ;
      RECT 0.261 0.486 0.345 0.522 ;
      RECT 0.345 0.486 0.364 0.522 ;
      RECT 0.364 0.486 0.597 0.522 ;
      RECT 0.597 0.486 0.639 0.522 ;
      RECT 0.639 0.486 0.726 0.522 ;
      RECT 0.726 0.486 0.912 0.522 ;
      RECT 0.912 0.486 0.977 0.522 ;
      RECT 0.977 0.486 1.099 0.522 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT -0.007 -0.018 1.099 0.018 ;
    END
  END VSS
  OBS
    LAYER MINT1 ;
      RECT 0.096 0.138 0.744 0.156 ;
      RECT 0.054 0.348 0.744 0.366 ;
    LAYER M1 ;
      RECT 0.117 0.047 0.135 0.457 ;
      RECT 0.201 0.047 0.219 0.457 ;
      RECT 0.285 0.080 0.303 0.098 ;
      RECT 0.285 0.098 0.303 0.240 ;
      RECT 0.285 0.240 0.303 0.440 ;
      RECT 0.303 0.080 0.537 0.098 ;
      RECT 0.537 0.080 0.555 0.098 ;
      RECT 0.537 0.098 0.555 0.240 ;
      RECT 0.621 0.180 0.639 0.377 ;
      RECT 0.705 0.127 0.726 0.213 ;
      RECT 0.705 0.258 0.726 0.390 ;
      RECT 0.831 0.122 0.849 0.209 ;
      RECT 0.789 0.259 0.807 0.377 ;
      RECT 0.789 0.377 0.807 0.395 ;
      RECT 0.807 0.377 0.957 0.395 ;
      RECT 0.957 0.047 0.975 0.087 ;
      RECT 0.957 0.087 0.975 0.259 ;
      RECT 0.957 0.259 0.975 0.377 ;
      RECT 0.957 0.377 0.975 0.395 ;
      RECT 0.975 0.087 0.977 0.259 ;
      RECT 0.975 0.259 0.977 0.377 ;
      RECT 0.975 0.377 0.977 0.395 ;
      RECT 0.030 0.054 0.032 0.091 ;
      RECT 0.030 0.091 0.032 0.116 ;
      RECT 0.032 0.054 0.052 0.091 ;
      RECT 0.032 0.091 0.052 0.116 ;
      RECT 0.032 0.372 0.052 0.398 ;
      RECT 0.032 0.398 0.052 0.450 ;
      RECT 0.052 0.054 0.054 0.091 ;
      RECT 0.052 0.091 0.054 0.116 ;
      RECT 0.052 0.372 0.054 0.398 ;
      RECT 0.054 0.091 0.075 0.116 ;
      RECT 0.054 0.372 0.075 0.398 ;
      RECT 0.075 0.091 0.093 0.116 ;
      RECT 0.075 0.116 0.093 0.372 ;
      RECT 0.075 0.372 0.093 0.398 ;
      RECT 0.243 0.127 0.261 0.324 ;
      RECT 0.327 0.264 0.345 0.387 ;
      RECT 0.345 0.127 0.364 0.200 ;
      RECT 0.495 0.169 0.513 0.240 ;
      RECT 0.399 0.180 0.417 0.377 ;
      RECT 0.399 0.377 0.417 0.395 ;
      RECT 0.417 0.377 0.576 0.395 ;
      RECT 0.576 0.377 0.579 0.395 ;
      RECT 0.576 0.395 0.579 0.450 ;
      RECT 0.579 0.063 0.597 0.180 ;
      RECT 0.579 0.180 0.597 0.377 ;
      RECT 0.579 0.377 0.597 0.395 ;
      RECT 0.579 0.395 0.597 0.450 ;
      RECT 0.663 0.075 0.681 0.093 ;
      RECT 0.663 0.093 0.681 0.240 ;
      RECT 0.663 0.240 0.681 0.441 ;
      RECT 0.681 0.075 0.887 0.093 ;
      RECT 0.887 0.075 0.906 0.093 ;
      RECT 0.887 0.093 0.906 0.240 ;
      RECT 0.726 0.419 0.912 0.437 ;
    LAYER V1 ;
      RECT 0.075 0.348 0.093 0.366 ;
      RECT 0.117 0.138 0.135 0.156 ;
      RECT 0.243 0.138 0.261 0.156 ;
      RECT 0.327 0.348 0.345 0.366 ;
      RECT 0.345 0.138 0.364 0.156 ;
      RECT 0.495 0.180 0.513 0.198 ;
      RECT 0.621 0.348 0.639 0.366 ;
      RECT 0.705 0.138 0.723 0.156 ;
      RECT 0.705 0.348 0.723 0.366 ;
      RECT 0.831 0.180 0.849 0.198 ;
  END
END DFFSNQ_X1

MACRO INV_X1
  CLASS core ;
  FOREIGN INV_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.126 BY 0.384 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.096 0.051 0.288   ; 
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.057 0.093 0.320   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.133 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.133 0.014   ; 
    END
  END VSS
END INV_X1

MACRO INV_X2
  CLASS core ;
  FOREIGN INV_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.126 BY 0.384 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.025 0.096 0.038 0.288   ; 
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.056 0.065 0.070 0.288   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.005 0.370 0.131 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.005 -0.014 0.131 0.014   ; 
    END
  END VSS
END INV_X2

MACRO INV_X4
  CLASS core ;
  FOREIGN INV_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.126 BY 0.384 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.016 0.128 0.026 0.184   ; 
RECT 0.016 0.184 0.026 0.198   ; 
RECT 0.016 0.198 0.026 0.256   ; 
RECT 0.026 0.184 0.078 0.198   ; 
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.013 0.071 0.019 0.100   ; 
RECT 0.019 0.071 0.100 0.100   ; 
RECT 0.019 0.284 0.100 0.313   ; 
RECT 0.100 0.071 0.110 0.100   ; 
RECT 0.100 0.100 0.110 0.284   ; 
RECT 0.100 0.284 0.110 0.313   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.003 0.370 0.129 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.003 -0.014 0.129 0.014   ; 
    END
  END VSS
END INV_X4

MACRO INV_X8
  CLASS core ;
  FOREIGN INV_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.126 BY 0.384 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.022 0.097 0.028 0.198   ; 
RECT 0.022 0.198 0.028 0.228   ; 
RECT 0.022 0.228 0.028 0.288   ; 
RECT 0.028 0.198 0.091 0.228   ; 
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.008 0.315 0.011 0.329   ; 
RECT 0.011 0.055 0.110 0.069   ; 
RECT 0.011 0.315 0.110 0.329   ; 
RECT 0.110 0.055 0.117 0.069   ; 
RECT 0.110 0.069 0.117 0.315   ; 
RECT 0.110 0.315 0.117 0.329   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 0.370 0.128 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 -0.014 0.128 0.014   ; 
    END
  END VSS
END INV_X8

MACRO INV_X12
  CLASS core ;
  FOREIGN INV_X12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.168 BY 0.384 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.021 0.096 0.027 0.184   ; 
RECT 0.021 0.184 0.027 0.198   ; 
RECT 0.021 0.198 0.027 0.288   ; 
RECT 0.027 0.184 0.129 0.198   ; 
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.010 0.051 0.152 0.065   ; 
RECT 0.010 0.318 0.152 0.334   ; 
RECT 0.152 0.051 0.160 0.065   ; 
RECT 0.152 0.065 0.160 0.318   ; 
RECT 0.152 0.318 0.160 0.334   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 0.370 0.170 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 -0.014 0.170 0.014   ; 
    END
  END VSS
END INV_X12

MACRO INV_X16
  CLASS core ;
  FOREIGN INV_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.168 BY 0.384 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.007 0.128 0.011 0.185   ; 
RECT 0.007 0.185 0.011 0.199   ; 
RECT 0.007 0.199 0.011 0.281   ; 
RECT 0.011 0.185 0.137 0.199   ; 
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.001 0.370 0.156 0.398   ; 
RECT 0.156 0.370 0.169 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.001 -0.014 0.169 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.008 0.050 0.151 0.066   ; 
RECT 0.008 0.311 0.151 0.341   ; 
RECT 0.151 0.050 0.156 0.066   ; 
RECT 0.151 0.066 0.156 0.311   ; 
RECT 0.151 0.311 0.156 0.341   ; 
      LAYER M1 ;
RECT 0.008 0.050 0.151 0.066   ; 
RECT 0.008 0.311 0.151 0.341   ; 
RECT 0.151 0.050 0.156 0.066   ; 
RECT 0.151 0.066 0.156 0.311   ; 
RECT 0.151 0.311 0.156 0.341   ; 
  END
END INV_X16

MACRO LHQ_X1
  CLASS core ;
  FOREIGN LHQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.588 BY 0.384 ; 
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.159 0.080 0.177 0.256   ; 
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
RECT 0.033 0.128 0.051 0.256   ; 
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.537 0.065 0.555 0.319   ; 
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.513 0.398   ; 
RECT 0.513 0.370 0.595 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.595 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.032 0.278 0.033 0.292   ; 
RECT 0.032 0.292 0.033 0.352   ; 
RECT 0.033 0.032 0.051 0.046   ; 
RECT 0.033 0.046 0.051 0.092   ; 
RECT 0.033 0.092 0.051 0.106   ; 
RECT 0.033 0.278 0.051 0.292   ; 
RECT 0.033 0.292 0.051 0.352   ; 
RECT 0.051 0.032 0.052 0.046   ; 
RECT 0.051 0.092 0.052 0.106   ; 
RECT 0.051 0.278 0.052 0.292   ; 
RECT 0.051 0.292 0.052 0.352   ; 
RECT 0.052 0.032 0.075 0.046   ; 
RECT 0.052 0.092 0.075 0.106   ; 
RECT 0.052 0.278 0.075 0.292   ; 
RECT 0.075 0.032 0.093 0.046   ; 
RECT 0.075 0.092 0.093 0.106   ; 
RECT 0.075 0.106 0.093 0.161   ; 
RECT 0.075 0.161 0.093 0.175   ; 
RECT 0.075 0.175 0.093 0.207   ; 
RECT 0.075 0.207 0.093 0.278   ; 
RECT 0.075 0.278 0.093 0.292   ; 
RECT 0.093 0.032 0.213 0.046   ; 
RECT 0.213 0.032 0.231 0.046   ; 
RECT 0.213 0.046 0.231 0.092   ; 
RECT 0.213 0.092 0.231 0.106   ; 
RECT 0.213 0.106 0.231 0.161   ; 
RECT 0.213 0.161 0.231 0.175   ; 
RECT 0.231 0.161 0.243 0.175   ; 
RECT 0.243 0.161 0.261 0.175   ; 
RECT 0.243 0.175 0.261 0.207   ; 
RECT 0.348 0.057 0.366 0.071   ; 
RECT 0.348 0.071 0.366 0.247   ; 
RECT 0.366 0.057 0.453 0.071   ; 
RECT 0.453 0.057 0.471 0.071   ; 
RECT 0.453 0.071 0.471 0.247   ; 
RECT 0.453 0.247 0.471 0.296   ; 
RECT 0.117 0.068 0.135 0.230   ; 
RECT 0.117 0.230 0.135 0.278   ; 
RECT 0.117 0.278 0.135 0.292   ; 
RECT 0.135 0.278 0.201 0.292   ; 
RECT 0.201 0.230 0.223 0.278   ; 
RECT 0.201 0.278 0.223 0.292   ; 
RECT 0.180 0.319 0.255 0.333   ; 
RECT 0.255 0.057 0.306 0.086   ; 
RECT 0.255 0.319 0.306 0.333   ; 
RECT 0.306 0.057 0.324 0.086   ; 
RECT 0.306 0.086 0.324 0.153   ; 
RECT 0.306 0.153 0.324 0.318   ; 
RECT 0.306 0.318 0.324 0.319   ; 
RECT 0.306 0.319 0.324 0.333   ; 
RECT 0.324 0.318 0.495 0.319   ; 
RECT 0.324 0.319 0.495 0.333   ; 
RECT 0.495 0.153 0.513 0.318   ; 
RECT 0.495 0.318 0.513 0.319   ; 
RECT 0.495 0.319 0.513 0.333   ; 
      LAYER M1 ;
RECT 0.032 0.278 0.033 0.292   ; 
RECT 0.032 0.292 0.033 0.352   ; 
RECT 0.033 0.032 0.051 0.046   ; 
RECT 0.033 0.046 0.051 0.092   ; 
RECT 0.033 0.092 0.051 0.106   ; 
RECT 0.033 0.278 0.051 0.292   ; 
RECT 0.033 0.292 0.051 0.352   ; 
RECT 0.051 0.032 0.052 0.046   ; 
RECT 0.051 0.092 0.052 0.106   ; 
RECT 0.051 0.278 0.052 0.292   ; 
RECT 0.051 0.292 0.052 0.352   ; 
RECT 0.052 0.032 0.075 0.046   ; 
RECT 0.052 0.092 0.075 0.106   ; 
RECT 0.052 0.278 0.075 0.292   ; 
RECT 0.075 0.032 0.093 0.046   ; 
RECT 0.075 0.092 0.093 0.106   ; 
RECT 0.075 0.106 0.093 0.161   ; 
RECT 0.075 0.161 0.093 0.175   ; 
RECT 0.075 0.175 0.093 0.207   ; 
RECT 0.075 0.207 0.093 0.278   ; 
RECT 0.075 0.278 0.093 0.292   ; 
RECT 0.093 0.032 0.213 0.046   ; 
RECT 0.213 0.032 0.231 0.046   ; 
RECT 0.213 0.046 0.231 0.092   ; 
RECT 0.213 0.092 0.231 0.106   ; 
RECT 0.213 0.106 0.231 0.161   ; 
RECT 0.213 0.161 0.231 0.175   ; 
RECT 0.231 0.161 0.243 0.175   ; 
RECT 0.243 0.161 0.261 0.175   ; 
RECT 0.243 0.175 0.261 0.207   ; 
RECT 0.348 0.057 0.366 0.071   ; 
RECT 0.348 0.071 0.366 0.247   ; 
RECT 0.366 0.057 0.453 0.071   ; 
RECT 0.453 0.057 0.471 0.071   ; 
RECT 0.453 0.071 0.471 0.247   ; 
RECT 0.453 0.247 0.471 0.296   ; 
RECT 0.117 0.068 0.135 0.230   ; 
RECT 0.117 0.230 0.135 0.278   ; 
RECT 0.117 0.278 0.135 0.292   ; 
RECT 0.135 0.278 0.201 0.292   ; 
RECT 0.201 0.230 0.223 0.278   ; 
RECT 0.201 0.278 0.223 0.292   ; 
RECT 0.180 0.319 0.255 0.333   ; 
RECT 0.255 0.057 0.306 0.086   ; 
RECT 0.255 0.319 0.306 0.333   ; 
RECT 0.306 0.057 0.324 0.086   ; 
RECT 0.306 0.086 0.324 0.153   ; 
RECT 0.306 0.153 0.324 0.318   ; 
RECT 0.306 0.318 0.324 0.319   ; 
RECT 0.306 0.319 0.324 0.333   ; 
RECT 0.324 0.318 0.495 0.319   ; 
RECT 0.324 0.319 0.495 0.333   ; 
RECT 0.495 0.153 0.513 0.318   ; 
RECT 0.495 0.318 0.513 0.319   ; 
RECT 0.495 0.319 0.513 0.333   ; 
  END
END LHQ_X1

MACRO MUX2_X1
  CLASS core ;
  FOREIGN MUX2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.546 BY 0.384 ;
  PIN I0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 0.373 0.121 0.395 0.263 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 0.085 0.128 0.107 0.224 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.121 0.036 0.329 ;
        RECT 0.018 0.329 0.036 0.343 ;
        RECT 0.036 0.329 0.146 0.343 ;
      LAYER V1 ;
        RECT 0.098 0.329 0.135 0.343 ;
      LAYER MINT1 ;
        RECT 0.077 0.408 0.259 0.432 ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT 0.469 0.096 0.491 0.319 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT -0.007 0.370 0.303 0.398 ;
      RECT 0.303 0.370 0.345 0.398 ;
      RECT 0.345 0.370 0.513 0.398 ;
      RECT 0.513 0.370 0.553 0.398 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT -0.007 -0.014 0.553 0.014 ;
    END
  END VSS
  OBS
    LAYER MINT1 ;
      RECT 0.180 0.222 0.366 0.240 ;
    LAYER M1 ;
      RECT 0.052 0.081 0.065 0.095 ;
      RECT 0.065 0.081 0.103 0.095 ;
      RECT 0.065 0.246 0.103 0.260 ;
      RECT 0.065 0.260 0.103 0.288 ;
      RECT 0.103 0.081 0.201 0.095 ;
      RECT 0.103 0.246 0.201 0.260 ;
      RECT 0.201 0.081 0.219 0.095 ;
      RECT 0.201 0.095 0.219 0.246 ;
      RECT 0.201 0.246 0.219 0.260 ;
      RECT 0.190 0.329 0.285 0.352 ;
      RECT 0.285 0.153 0.303 0.329 ;
      RECT 0.285 0.329 0.303 0.352 ;
      RECT 0.327 0.137 0.345 0.214 ;
      RECT 0.243 0.043 0.261 0.073 ;
      RECT 0.243 0.073 0.261 0.247 ;
      RECT 0.243 0.247 0.261 0.307 ;
      RECT 0.261 0.043 0.495 0.073 ;
      RECT 0.495 0.043 0.513 0.073 ;
      RECT 0.495 0.073 0.513 0.247 ;
    LAYER V1 ;
      RECT 0.201 0.169 0.219 0.183 ;
      RECT 0.201 0.329 0.238 0.343 ;
      RECT 0.327 0.169 0.345 0.183 ;
  END
END MUX2_X1

MACRO NAND2_X1
  CLASS core ;
  FOREIGN NAND2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.168 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.128 0.135 0.287   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.128 0.051 0.287   ; 
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.067 0.093 0.096   ; 
RECT 0.075 0.096 0.093 0.319   ; 
RECT 0.093 0.067 0.116 0.096   ; 
RECT 0.116 0.032 0.137 0.067   ; 
RECT 0.116 0.067 0.137 0.096   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.175 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.175 0.014   ; 
    END
  END VSS
END NAND2_X1

MACRO NAND2_X2
  CLASS core ;
  FOREIGN NAND2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.168 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.078 0.113 0.090 0.277   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.022 0.137 0.034 0.338   ; 
RECT 0.022 0.338 0.034 0.352   ; 
RECT 0.034 0.338 0.134 0.352   ; 
RECT 0.134 0.137 0.146 0.338   ; 
RECT 0.134 0.338 0.146 0.352   ; 
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.050 0.062 0.062 0.091   ; 
RECT 0.050 0.091 0.062 0.212   ; 
RECT 0.050 0.212 0.062 0.299   ; 
RECT 0.050 0.299 0.062 0.320   ; 
RECT 0.062 0.062 0.106 0.091   ; 
RECT 0.062 0.299 0.106 0.320   ; 
RECT 0.106 0.062 0.118 0.091   ; 
RECT 0.106 0.212 0.118 0.299   ; 
RECT 0.106 0.299 0.118 0.320   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.370 0.172 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.014 0.172 0.014   ; 
    END
  END VSS
END NAND2_X2

MACRO NAND3_X1
  CLASS core ;
  FOREIGN NAND3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.159 0.160 0.177 0.224   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.128 0.135 0.256   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.108 0.051 0.287   ; 
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.041 0.093 0.055   ; 
RECT 0.075 0.055 0.093 0.128   ; 
RECT 0.075 0.128 0.093 0.256   ; 
RECT 0.075 0.256 0.093 0.338   ; 
RECT 0.075 0.338 0.093 0.352   ; 
RECT 0.093 0.041 0.159 0.055   ; 
RECT 0.093 0.338 0.159 0.352   ; 
RECT 0.159 0.032 0.200 0.041   ; 
RECT 0.159 0.041 0.200 0.055   ; 
RECT 0.159 0.338 0.200 0.352   ; 
RECT 0.200 0.032 0.201 0.041   ; 
RECT 0.200 0.041 0.201 0.055   ; 
RECT 0.200 0.055 0.201 0.128   ; 
RECT 0.200 0.338 0.201 0.352   ; 
RECT 0.201 0.032 0.219 0.041   ; 
RECT 0.201 0.041 0.219 0.055   ; 
RECT 0.201 0.055 0.219 0.128   ; 
RECT 0.201 0.256 0.219 0.338   ; 
RECT 0.201 0.338 0.219 0.352   ; 
RECT 0.219 0.032 0.221 0.041   ; 
RECT 0.219 0.041 0.221 0.055   ; 
RECT 0.219 0.055 0.221 0.128   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.259 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.259 0.014   ; 
    END
  END VSS
END NAND3_X1

MACRO NAND3_X2
  CLASS core ;
  FOREIGN NAND3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.218 0.160 0.230 0.256   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.132 0.124 0.148 0.256   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.050 0.128 0.062 0.256   ; 
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.012 0.284 0.160 0.313   ; 
RECT 0.160 0.284 0.190 0.313   ; 
RECT 0.190 0.093 0.202 0.284   ; 
RECT 0.190 0.284 0.202 0.313   ; 
RECT 0.202 0.284 0.216 0.313   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.370 0.160 0.398   ; 
RECT 0.160 0.370 0.230 0.398   ; 
RECT 0.230 0.370 0.256 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.014 0.256 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.092 0.056 0.218 0.070   ; 
RECT 0.218 0.056 0.230 0.070   ; 
RECT 0.218 0.070 0.230 0.113   ; 
RECT 0.022 0.088 0.160 0.104   ; 
      LAYER M1 ;
RECT 0.092 0.056 0.218 0.070   ; 
RECT 0.218 0.056 0.230 0.070   ; 
RECT 0.218 0.070 0.230 0.113   ; 
RECT 0.022 0.088 0.160 0.104   ; 
  END
END NAND3_X2

MACRO NAND4_X1
  CLASS core ;
  FOREIGN NAND4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.243 0.128 0.261 0.287   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.159 0.121 0.177 0.256   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.097 0.135 0.224   ; 
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.097 0.051 0.287   ; 
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.256 0.093 0.322   ; 
RECT 0.075 0.322 0.093 0.352   ; 
RECT 0.093 0.322 0.201 0.352   ; 
RECT 0.201 0.082 0.219 0.096   ; 
RECT 0.201 0.096 0.219 0.256   ; 
RECT 0.201 0.256 0.219 0.322   ; 
RECT 0.201 0.322 0.219 0.352   ; 
RECT 0.219 0.082 0.240 0.096   ; 
RECT 0.240 0.032 0.264 0.082   ; 
RECT 0.240 0.082 0.264 0.096   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.301 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.301 0.014   ; 
    END
  END VSS
END NAND4_X1

MACRO NAND4_X2
  CLASS core ;
  FOREIGN NAND4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.233 0.179 0.248 0.256   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.155 0.170 0.166 0.263   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.074 0.121 0.086 0.256   ; 
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.021 0.129 0.033 0.256   ; 
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.047 0.277 0.060 0.288   ; 
RECT 0.047 0.288 0.060 0.319   ; 
RECT 0.047 0.319 0.060 0.333   ; 
RECT 0.060 0.319 0.181 0.333   ; 
RECT 0.181 0.147 0.193 0.161   ; 
RECT 0.181 0.161 0.193 0.274   ; 
RECT 0.181 0.274 0.193 0.277   ; 
RECT 0.181 0.277 0.193 0.288   ; 
RECT 0.181 0.319 0.193 0.333   ; 
RECT 0.193 0.147 0.235 0.161   ; 
RECT 0.193 0.274 0.235 0.277   ; 
RECT 0.193 0.277 0.235 0.288   ; 
RECT 0.193 0.319 0.235 0.333   ; 
RECT 0.235 0.147 0.246 0.161   ; 
RECT 0.235 0.274 0.246 0.277   ; 
RECT 0.235 0.277 0.246 0.288   ; 
RECT 0.235 0.288 0.246 0.319   ; 
RECT 0.235 0.319 0.246 0.333   ; 
RECT 0.246 0.147 0.273 0.161   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.370 0.274 0.398   ; 
RECT 0.274 0.370 0.298 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.014 0.298 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.020 0.051 0.033 0.065   ; 
RECT 0.020 0.065 0.033 0.107   ; 
RECT 0.033 0.051 0.180 0.065   ; 
RECT 0.114 0.115 0.261 0.129   ; 
RECT 0.261 0.032 0.274 0.115   ; 
RECT 0.261 0.115 0.274 0.129   ; 
RECT 0.061 0.083 0.206 0.097   ; 
      LAYER M1 ;
RECT 0.020 0.051 0.033 0.065   ; 
RECT 0.020 0.065 0.033 0.107   ; 
RECT 0.033 0.051 0.180 0.065   ; 
RECT 0.114 0.115 0.261 0.129   ; 
RECT 0.261 0.032 0.274 0.115   ; 
RECT 0.261 0.115 0.274 0.129   ; 
RECT 0.061 0.083 0.206 0.097   ; 
  END
END NAND4_X2

MACRO NOR2_X1
  CLASS core ;
  FOREIGN NOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.168 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.097 0.135 0.256   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.097 0.051 0.256   ; 
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.065 0.093 0.288   ; 
RECT 0.075 0.288 0.093 0.318   ; 
RECT 0.093 0.288 0.116 0.318   ; 
RECT 0.116 0.288 0.137 0.318   ; 
RECT 0.116 0.318 0.137 0.352   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.175 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.175 0.014   ; 
    END
  END VSS
END NOR2_X1

MACRO NOR2_X2
  CLASS core ;
  FOREIGN NOR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.168 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.078 0.107 0.090 0.256   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.022 0.032 0.034 0.046   ; 
RECT 0.022 0.046 0.034 0.247   ; 
RECT 0.034 0.032 0.134 0.046   ; 
RECT 0.134 0.032 0.146 0.046   ; 
RECT 0.134 0.046 0.146 0.247   ; 
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.050 0.064 0.062 0.078   ; 
RECT 0.050 0.078 0.062 0.172   ; 
RECT 0.050 0.172 0.062 0.278   ; 
RECT 0.050 0.278 0.062 0.292   ; 
RECT 0.062 0.064 0.077 0.078   ; 
RECT 0.062 0.278 0.077 0.292   ; 
RECT 0.077 0.064 0.091 0.078   ; 
RECT 0.077 0.278 0.091 0.292   ; 
RECT 0.077 0.292 0.091 0.320   ; 
RECT 0.091 0.064 0.106 0.078   ; 
RECT 0.106 0.064 0.118 0.078   ; 
RECT 0.106 0.078 0.118 0.172   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.370 0.172 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.014 0.172 0.014   ; 
    END
  END VSS
END NOR2_X2

MACRO NOR3_X1
  CLASS core ;
  FOREIGN NOR3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.159 0.160 0.177 0.224   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.097 0.135 0.276   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.097 0.051 0.276   ; 
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.032 0.093 0.046   ; 
RECT 0.075 0.046 0.093 0.128   ; 
RECT 0.075 0.128 0.093 0.256   ; 
RECT 0.075 0.256 0.093 0.307   ; 
RECT 0.075 0.307 0.093 0.321   ; 
RECT 0.093 0.032 0.199 0.046   ; 
RECT 0.093 0.307 0.199 0.321   ; 
RECT 0.199 0.032 0.200 0.046   ; 
RECT 0.199 0.046 0.200 0.128   ; 
RECT 0.199 0.307 0.200 0.321   ; 
RECT 0.200 0.032 0.221 0.046   ; 
RECT 0.200 0.046 0.221 0.128   ; 
RECT 0.200 0.256 0.221 0.307   ; 
RECT 0.200 0.307 0.221 0.321   ; 
RECT 0.200 0.321 0.221 0.352   ; 
RECT 0.221 0.032 0.221 0.046   ; 
RECT 0.221 0.046 0.221 0.128   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.259 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.259 0.014   ; 
    END
  END VSS
END NOR3_X1

MACRO NOR3_X2
  CLASS core ;
  FOREIGN NOR3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.218 0.128 0.230 0.224   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.134 0.128 0.146 0.257   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.022 0.128 0.034 0.260   ; 
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.038 0.077 0.190 0.106   ; 
RECT 0.190 0.077 0.202 0.106   ; 
RECT 0.190 0.106 0.202 0.288   ; 
RECT 0.202 0.077 0.214 0.106   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.370 0.230 0.398   ; 
RECT 0.230 0.370 0.256 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.014 0.256 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.092 0.313 0.218 0.328   ; 
RECT 0.218 0.258 0.230 0.313   ; 
RECT 0.218 0.313 0.230 0.328   ; 
RECT 0.038 0.279 0.166 0.296   ; 
      LAYER M1 ;
RECT 0.092 0.313 0.218 0.328   ; 
RECT 0.218 0.258 0.230 0.313   ; 
RECT 0.218 0.313 0.230 0.328   ; 
RECT 0.038 0.279 0.166 0.296   ; 
  END
END NOR3_X2

MACRO NOR4_X1
  CLASS core ;
  FOREIGN NOR4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.243 0.097 0.261 0.256   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.159 0.097 0.177 0.256   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.128 0.135 0.287   ; 
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.097 0.051 0.287   ; 
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.032 0.093 0.051   ; 
RECT 0.075 0.051 0.093 0.108   ; 
RECT 0.093 0.032 0.201 0.051   ; 
RECT 0.201 0.032 0.219 0.051   ; 
RECT 0.201 0.051 0.219 0.108   ; 
RECT 0.201 0.108 0.219 0.288   ; 
RECT 0.201 0.288 0.219 0.302   ; 
RECT 0.219 0.288 0.240 0.302   ; 
RECT 0.240 0.288 0.264 0.302   ; 
RECT 0.240 0.302 0.264 0.352   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.301 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.301 0.014   ; 
    END
  END VSS
END NOR4_X1

MACRO NOR4_X2
  CLASS core ;
  FOREIGN NOR4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.233 0.128 0.248 0.203   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.155 0.121 0.166 0.219   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.101 0.121 0.113 0.263   ; 
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.074 0.128 0.086 0.258   ; 
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.047 0.051 0.060 0.065   ; 
RECT 0.047 0.065 0.060 0.096   ; 
RECT 0.047 0.096 0.060 0.107   ; 
RECT 0.060 0.051 0.181 0.065   ; 
RECT 0.181 0.051 0.193 0.065   ; 
RECT 0.181 0.096 0.193 0.107   ; 
RECT 0.181 0.107 0.193 0.110   ; 
RECT 0.181 0.110 0.193 0.221   ; 
RECT 0.181 0.221 0.193 0.235   ; 
RECT 0.193 0.051 0.235 0.065   ; 
RECT 0.193 0.096 0.235 0.107   ; 
RECT 0.193 0.107 0.235 0.110   ; 
RECT 0.193 0.221 0.235 0.235   ; 
RECT 0.235 0.051 0.246 0.065   ; 
RECT 0.235 0.065 0.246 0.096   ; 
RECT 0.235 0.096 0.246 0.107   ; 
RECT 0.235 0.107 0.246 0.110   ; 
RECT 0.235 0.221 0.246 0.235   ; 
RECT 0.246 0.221 0.277 0.235   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.370 0.180 0.398   ; 
RECT 0.180 0.370 0.206 0.398   ; 
RECT 0.206 0.370 0.274 0.398   ; 
RECT 0.274 0.370 0.298 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.014 0.298 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.088 0.285 0.206 0.301   ; 
RECT 0.020 0.277 0.033 0.319   ; 
RECT 0.020 0.319 0.033 0.333   ; 
RECT 0.033 0.319 0.180 0.333   ; 
RECT 0.141 0.253 0.261 0.267   ; 
RECT 0.261 0.253 0.274 0.267   ; 
RECT 0.261 0.267 0.274 0.343   ; 
      LAYER M1 ;
RECT 0.088 0.285 0.206 0.301   ; 
RECT 0.020 0.277 0.033 0.319   ; 
RECT 0.020 0.319 0.033 0.333   ; 
RECT 0.033 0.319 0.180 0.333   ; 
RECT 0.141 0.253 0.261 0.267   ; 
RECT 0.261 0.253 0.274 0.267   ; 
RECT 0.261 0.267 0.274 0.343   ; 
  END
END NOR4_X2


MACRO OAI21_X1
  CLASS core ;
  FOREIGN OAI21_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.128 0.135 0.288   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.128 0.051 0.317   ; 
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.201 0.128 0.219 0.288   ; 
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.128 0.093 0.318   ; 
RECT 0.075 0.318 0.093 0.334   ; 
RECT 0.093 0.318 0.196 0.334   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.196 0.398   ; 
RECT 0.196 0.370 0.259 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.259 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.033 0.036 0.051 0.078   ; 
RECT 0.033 0.078 0.051 0.094   ; 
RECT 0.051 0.078 0.196 0.094   ; 
      LAYER M1 ;
RECT 0.033 0.036 0.051 0.078   ; 
RECT 0.033 0.078 0.051 0.094   ; 
RECT 0.051 0.078 0.196 0.094   ; 
  END
END OAI21_X1

MACRO OAI21_X2
  CLASS core ;
  FOREIGN OAI21_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.160 0.160 0.176 0.224   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.106 0.121 0.118 0.142   ; 
RECT 0.106 0.142 0.118 0.251   ; 
RECT 0.106 0.251 0.118 0.265   ; 
RECT 0.118 0.251 0.218 0.265   ; 
RECT 0.218 0.142 0.230 0.251   ; 
RECT 0.218 0.251 0.230 0.265   ; 
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.050 0.128 0.062 0.263   ; 
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.013 0.285 0.078 0.301   ; 
RECT 0.078 0.083 0.090 0.097   ; 
RECT 0.078 0.097 0.090 0.139   ; 
RECT 0.078 0.139 0.090 0.285   ; 
RECT 0.078 0.285 0.090 0.301   ; 
RECT 0.090 0.083 0.186 0.097   ; 
RECT 0.090 0.285 0.186 0.301   ; 
RECT 0.186 0.083 0.190 0.097   ; 
RECT 0.190 0.083 0.202 0.097   ; 
RECT 0.190 0.097 0.202 0.139   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.370 0.234 0.398   ; 
RECT 0.234 0.370 0.256 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.014 0.256 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.021 0.051 0.035 0.065   ; 
RECT 0.021 0.065 0.035 0.107   ; 
RECT 0.035 0.051 0.218 0.065   ; 
RECT 0.218 0.051 0.230 0.065   ; 
RECT 0.218 0.065 0.230 0.107   ; 
RECT 0.218 0.107 0.230 0.107   ; 
RECT 0.064 0.319 0.234 0.333   ; 
      LAYER M1 ;
RECT 0.021 0.051 0.035 0.065   ; 
RECT 0.021 0.065 0.035 0.107   ; 
RECT 0.035 0.051 0.218 0.065   ; 
RECT 0.218 0.051 0.230 0.065   ; 
RECT 0.218 0.065 0.230 0.107   ; 
RECT 0.218 0.107 0.230 0.107   ; 
RECT 0.064 0.319 0.234 0.333   ; 
  END
END OAI21_X2

MACRO OAI22_X1
  CLASS core ;
  FOREIGN OAI22_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.159 0.100 0.177 0.288   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.243 0.140 0.261 0.288   ; 
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.096 0.135 0.256   ; 
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.032 0.096 0.052 0.288   ; 
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.092 0.319 0.201 0.333   ; 
RECT 0.201 0.091 0.219 0.319   ; 
RECT 0.201 0.319 0.219 0.333   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.261 0.398   ; 
RECT 0.261 0.370 0.301 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.301 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.033 0.050 0.243 0.065   ; 
RECT 0.243 0.050 0.261 0.065   ; 
RECT 0.243 0.065 0.261 0.106   ; 
      LAYER M1 ;
RECT 0.033 0.050 0.243 0.065   ; 
RECT 0.243 0.050 0.261 0.065   ; 
RECT 0.243 0.065 0.261 0.106   ; 
  END
END OAI22_X1

MACRO OAI22_X2
  CLASS core ;
  FOREIGN OAI22_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.166 0.128 0.177 0.139   ; 
RECT 0.166 0.139 0.177 0.233   ; 
RECT 0.166 0.233 0.177 0.247   ; 
RECT 0.177 0.233 0.264 0.247   ; 
RECT 0.264 0.139 0.275 0.233   ; 
RECT 0.264 0.233 0.275 0.247   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.215 0.128 0.226 0.199   ; 
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.121 0.128 0.243   ; 
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.044 0.121 0.054 0.256   ; 
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.093 0.193 0.103 0.265   ; 
RECT 0.093 0.265 0.103 0.279   ; 
RECT 0.103 0.265 0.142 0.279   ; 
RECT 0.142 0.085 0.152 0.098   ; 
RECT 0.142 0.098 0.152 0.139   ; 
RECT 0.142 0.139 0.152 0.193   ; 
RECT 0.142 0.193 0.152 0.265   ; 
RECT 0.142 0.265 0.152 0.279   ; 
RECT 0.152 0.085 0.240 0.098   ; 
RECT 0.152 0.265 0.240 0.279   ; 
RECT 0.240 0.085 0.250 0.098   ; 
RECT 0.240 0.098 0.250 0.139   ; 
RECT 0.240 0.265 0.250 0.279   ; 
RECT 0.250 0.265 0.264 0.279   ; 
RECT 0.264 0.265 0.275 0.279   ; 
RECT 0.264 0.279 0.275 0.336   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.370 0.139 0.398   ; 
RECT 0.139 0.370 0.250 0.398   ; 
RECT 0.250 0.370 0.275 0.398   ; 
RECT 0.275 0.370 0.298 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.014 0.298 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.154 0.302 0.240 0.318   ; 
RECT 0.240 0.302 0.250 0.318   ; 
RECT 0.240 0.318 0.250 0.348   ; 
RECT 0.016 0.050 0.264 0.066   ; 
RECT 0.264 0.050 0.275 0.066   ; 
RECT 0.264 0.066 0.275 0.105   ; 
RECT 0.019 0.306 0.139 0.335   ; 
      LAYER M1 ;
RECT 0.154 0.302 0.240 0.318   ; 
RECT 0.240 0.302 0.250 0.318   ; 
RECT 0.240 0.318 0.250 0.348   ; 
RECT 0.016 0.050 0.264 0.066   ; 
RECT 0.264 0.050 0.275 0.066   ; 
RECT 0.264 0.066 0.275 0.105   ; 
RECT 0.019 0.306 0.139 0.335   ; 
  END
END OAI22_X2

MACRO OR2_X1
  CLASS core ;
  FOREIGN OR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.048 0.135 0.256   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.122 0.051 0.320   ; 
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.201 0.057 0.219 0.320   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.177 0.398   ; 
RECT 0.177 0.370 0.259 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.259 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.075 0.065 0.093 0.168   ; 
RECT 0.075 0.168 0.093 0.278   ; 
RECT 0.075 0.278 0.093 0.292   ; 
RECT 0.093 0.278 0.159 0.292   ; 
RECT 0.159 0.168 0.177 0.278   ; 
RECT 0.159 0.278 0.177 0.292   ; 
      LAYER M1 ;
RECT 0.075 0.065 0.093 0.168   ; 
RECT 0.075 0.168 0.093 0.278   ; 
RECT 0.075 0.278 0.093 0.292   ; 
RECT 0.093 0.278 0.159 0.292   ; 
RECT 0.159 0.168 0.177 0.278   ; 
RECT 0.159 0.278 0.177 0.292   ; 
  END
END OR2_X1

MACRO OR2_X2
  CLASS core ;
  FOREIGN OR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.064 0.121 0.080 0.256   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.028 0.128 0.044 0.256   ; 
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.170 0.032 0.172 0.068   ; 
RECT 0.170 0.319 0.172 0.352   ; 
RECT 0.172 0.032 0.188 0.068   ; 
RECT 0.172 0.068 0.188 0.319   ; 
RECT 0.172 0.319 0.188 0.352   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.006 0.370 0.152 0.398   ; 
RECT 0.152 0.370 0.258 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.006 -0.014 0.258 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.043 0.077 0.082 0.094   ; 
RECT 0.082 0.077 0.136 0.094   ; 
RECT 0.082 0.290 0.136 0.304   ; 
RECT 0.136 0.077 0.152 0.094   ; 
RECT 0.136 0.094 0.152 0.290   ; 
RECT 0.136 0.290 0.152 0.304   ; 
      LAYER M1 ;
RECT 0.043 0.077 0.082 0.094   ; 
RECT 0.082 0.077 0.136 0.094   ; 
RECT 0.082 0.290 0.136 0.304   ; 
RECT 0.136 0.077 0.152 0.094   ; 
RECT 0.136 0.094 0.152 0.290   ; 
RECT 0.136 0.290 0.152 0.304   ; 
  END
END OR2_X2

MACRO OR3_X1
  CLASS core ;
  FOREIGN OR3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.336 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.201 0.096 0.219 0.288   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.116 0.096 0.137 0.288   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.030 0.096 0.054 0.288   ; 
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.285 0.057 0.303 0.327   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.154 0.398   ; 
RECT 0.154 0.370 0.261 0.398   ; 
RECT 0.261 0.370 0.343 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.343 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.035 0.055 0.182 0.068   ; 
RECT 0.182 0.055 0.243 0.068   ; 
RECT 0.182 0.316 0.243 0.336   ; 
RECT 0.243 0.055 0.261 0.068   ; 
RECT 0.243 0.068 0.261 0.316   ; 
RECT 0.243 0.316 0.261 0.336   ; 
RECT 0.056 0.318 0.154 0.334   ; 
      LAYER M1 ;
RECT 0.035 0.055 0.182 0.068   ; 
RECT 0.182 0.055 0.243 0.068   ; 
RECT 0.182 0.316 0.243 0.336   ; 
RECT 0.243 0.055 0.261 0.068   ; 
RECT 0.243 0.068 0.261 0.316   ; 
RECT 0.243 0.316 0.261 0.336   ; 
RECT 0.056 0.318 0.154 0.334   ; 
  END
END OR3_X1

MACRO OR3_X2
  CLASS core ;
  FOREIGN OR3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.336 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.128 0.093 0.224   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.128 0.051 0.263   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.159 0.116 0.177 0.224   ; 
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.240 0.032 0.243 0.065   ; 
RECT 0.240 0.318 0.243 0.352   ; 
RECT 0.243 0.032 0.261 0.065   ; 
RECT 0.243 0.065 0.261 0.318   ; 
RECT 0.243 0.318 0.261 0.352   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.198 0.398   ; 
RECT 0.198 0.370 0.219 0.398   ; 
RECT 0.219 0.370 0.343 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.343 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.033 0.286 0.051 0.302   ; 
RECT 0.033 0.302 0.051 0.343   ; 
RECT 0.051 0.286 0.198 0.302   ; 
RECT 0.039 0.078 0.092 0.094   ; 
RECT 0.092 0.078 0.201 0.094   ; 
RECT 0.092 0.252 0.201 0.268   ; 
RECT 0.201 0.078 0.219 0.094   ; 
RECT 0.201 0.094 0.219 0.252   ; 
RECT 0.201 0.252 0.219 0.268   ; 
      LAYER M1 ;
RECT 0.033 0.286 0.051 0.302   ; 
RECT 0.033 0.302 0.051 0.343   ; 
RECT 0.051 0.286 0.198 0.302   ; 
RECT 0.039 0.078 0.092 0.094   ; 
RECT 0.092 0.078 0.201 0.094   ; 
RECT 0.092 0.252 0.201 0.268   ; 
RECT 0.201 0.078 0.219 0.094   ; 
RECT 0.201 0.094 0.219 0.252   ; 
RECT 0.201 0.252 0.219 0.268   ; 
  END
END OR3_X2

MACRO OR4_X1
  CLASS core ;
  FOREIGN OR4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.378 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.243 0.096 0.261 0.288   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.158 0.096 0.178 0.288   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.099 0.093 0.288   ; 
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.096 0.051 0.288   ; 
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.327 0.057 0.345 0.320   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.196 0.398   ; 
RECT 0.196 0.370 0.303 0.398   ; 
RECT 0.303 0.370 0.385 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.385 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.035 0.051 0.222 0.065   ; 
RECT 0.222 0.051 0.285 0.065   ; 
RECT 0.222 0.315 0.285 0.331   ; 
RECT 0.285 0.051 0.303 0.065   ; 
RECT 0.285 0.065 0.303 0.315   ; 
RECT 0.285 0.315 0.303 0.331   ; 
RECT 0.096 0.308 0.196 0.328   ; 
      LAYER M1 ;
RECT 0.035 0.051 0.222 0.065   ; 
RECT 0.222 0.051 0.285 0.065   ; 
RECT 0.222 0.315 0.285 0.331   ; 
RECT 0.285 0.051 0.303 0.065   ; 
RECT 0.285 0.065 0.303 0.315   ; 
RECT 0.285 0.315 0.303 0.331   ; 
RECT 0.096 0.308 0.196 0.328   ; 
  END
END OR4_X1

MACRO OR4_X2
  CLASS core ;
  FOREIGN OR4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.378 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.181 0.096 0.197 0.265   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.143 0.107 0.159 0.288   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.067 0.107 0.084 0.288   ; 
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.030 0.095 0.046 0.288   ; 
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.293 0.064 0.312 0.352   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.006 0.370 0.178 0.398   ; 
RECT 0.178 0.370 0.272 0.398   ; 
RECT 0.272 0.370 0.384 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.006 -0.014 0.384 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.086 0.312 0.178 0.341   ; 
RECT 0.032 0.043 0.202 0.072   ; 
RECT 0.202 0.043 0.255 0.072   ; 
RECT 0.202 0.284 0.255 0.312   ; 
RECT 0.255 0.043 0.272 0.072   ; 
RECT 0.255 0.072 0.272 0.284   ; 
RECT 0.255 0.284 0.272 0.312   ; 
      LAYER M1 ;
RECT 0.086 0.312 0.178 0.341   ; 
RECT 0.032 0.043 0.202 0.072   ; 
RECT 0.202 0.043 0.255 0.072   ; 
RECT 0.202 0.284 0.255 0.312   ; 
RECT 0.255 0.043 0.272 0.072   ; 
RECT 0.255 0.072 0.272 0.284   ; 
RECT 0.255 0.284 0.272 0.312   ; 
  END
END OR4_X2



MACRO TIEH
  CLASS core ;
  FOREIGN TIEH 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.126 BY 0.384 ; 
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.072 0.236 0.093 0.352   ; 
RECT 0.093 0.236 0.096 0.352   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.093 0.398   ; 
RECT 0.093 0.370 0.133 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.133 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.075 0.048 0.093 0.214   ; 
      LAYER M1 ;
RECT 0.075 0.048 0.093 0.214   ; 
  END
END TIEH

MACRO TIEL
  CLASS core ;
  FOREIGN TIEL 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.126 BY 0.384 ; 
  PIN Z
    DIRECTION INOUT ;
    PORT
      LAYER M1 ;
RECT 0.072 0.032 0.096 0.133   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.093 0.398   ; 
RECT 0.093 0.370 0.133 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.133 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.075 0.168 0.093 0.336   ; 
      LAYER M1 ;
RECT 0.075 0.168 0.093 0.336   ; 
  END
END TIEL

MACRO XNOR2_X1
  CLASS core ;
  FOREIGN XNOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.378 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.126 0.138 0.140   ; 
RECT 0.117 0.140 0.138 0.214   ; 
RECT 0.138 0.126 0.243 0.140   ; 
RECT 0.243 0.126 0.261 0.140   ; 
RECT 0.243 0.140 0.261 0.214   ; 
RECT 0.243 0.214 0.261 0.224   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.121 0.051 0.160   ; 
RECT 0.033 0.160 0.051 0.338   ; 
RECT 0.033 0.338 0.051 0.352   ; 
RECT 0.051 0.338 0.180 0.352   ; 
RECT 0.180 0.338 0.327 0.352   ; 
RECT 0.327 0.160 0.345 0.338   ; 
RECT 0.327 0.338 0.345 0.352   ; 
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.182 0.273 0.198 0.274   ; 
RECT 0.182 0.274 0.198 0.300   ; 
RECT 0.182 0.300 0.198 0.301   ; 
RECT 0.198 0.083 0.219 0.097   ; 
RECT 0.198 0.273 0.219 0.274   ; 
RECT 0.198 0.274 0.219 0.300   ; 
RECT 0.198 0.300 0.219 0.301   ; 
RECT 0.219 0.083 0.285 0.097   ; 
RECT 0.219 0.274 0.285 0.300   ; 
RECT 0.285 0.083 0.303 0.097   ; 
RECT 0.285 0.124 0.303 0.138   ; 
RECT 0.285 0.138 0.303 0.273   ; 
RECT 0.285 0.273 0.303 0.274   ; 
RECT 0.285 0.274 0.303 0.300   ; 
RECT 0.303 0.083 0.324 0.097   ; 
RECT 0.303 0.124 0.324 0.138   ; 
RECT 0.324 0.083 0.348 0.097   ; 
RECT 0.324 0.097 0.348 0.124   ; 
RECT 0.324 0.124 0.348 0.138   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.180 0.398   ; 
RECT 0.180 0.370 0.351 0.398   ; 
RECT 0.351 0.370 0.385 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.385 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.138 0.051 0.351 0.065   ; 
RECT 0.075 0.092 0.093 0.108   ; 
RECT 0.075 0.108 0.093 0.170   ; 
RECT 0.075 0.170 0.093 0.232   ; 
RECT 0.075 0.232 0.093 0.246   ; 
RECT 0.075 0.246 0.093 0.276   ; 
RECT 0.093 0.092 0.154 0.108   ; 
RECT 0.093 0.232 0.154 0.246   ; 
RECT 0.154 0.232 0.161 0.246   ; 
RECT 0.161 0.170 0.180 0.232   ; 
RECT 0.161 0.232 0.180 0.246   ; 
      LAYER M1 ;
RECT 0.138 0.051 0.351 0.065   ; 
RECT 0.075 0.092 0.093 0.108   ; 
RECT 0.075 0.108 0.093 0.170   ; 
RECT 0.075 0.170 0.093 0.232   ; 
RECT 0.075 0.232 0.093 0.246   ; 
RECT 0.075 0.246 0.093 0.276   ; 
RECT 0.093 0.092 0.154 0.108   ; 
RECT 0.093 0.232 0.154 0.246   ; 
RECT 0.154 0.232 0.161 0.246   ; 
RECT 0.161 0.170 0.180 0.232   ; 
RECT 0.161 0.232 0.180 0.246   ; 
  END
END XNOR2_X1

MACRO XOR2_X1
  CLASS core ;
  FOREIGN XOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.378 BY 0.384 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.172 0.138 0.243   ; 
RECT 0.117 0.243 0.138 0.257   ; 
RECT 0.138 0.243 0.180 0.257   ; 
RECT 0.180 0.243 0.243 0.257   ; 
RECT 0.243 0.160 0.261 0.172   ; 
RECT 0.243 0.172 0.261 0.243   ; 
RECT 0.243 0.243 0.261 0.257   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.032 0.051 0.046   ; 
RECT 0.033 0.046 0.051 0.224   ; 
RECT 0.033 0.224 0.051 0.263   ; 
RECT 0.051 0.032 0.327 0.046   ; 
RECT 0.327 0.032 0.345 0.046   ; 
RECT 0.327 0.046 0.345 0.224   ; 
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.180 0.082 0.207 0.082   ; 
RECT 0.180 0.082 0.207 0.111   ; 
RECT 0.207 0.082 0.219 0.082   ; 
RECT 0.207 0.082 0.219 0.111   ; 
RECT 0.207 0.287 0.219 0.301   ; 
RECT 0.219 0.082 0.285 0.111   ; 
RECT 0.219 0.287 0.285 0.301   ; 
RECT 0.285 0.082 0.303 0.111   ; 
RECT 0.285 0.111 0.303 0.246   ; 
RECT 0.285 0.246 0.303 0.260   ; 
RECT 0.285 0.287 0.303 0.301   ; 
RECT 0.303 0.246 0.326 0.260   ; 
RECT 0.303 0.287 0.326 0.301   ; 
RECT 0.326 0.246 0.346 0.260   ; 
RECT 0.326 0.260 0.346 0.287   ; 
RECT 0.326 0.287 0.346 0.301   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.370 0.351 0.398   ; 
RECT 0.351 0.370 0.385 0.398   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.014 0.385 0.014   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.161 0.319 0.351 0.333   ; 
RECT 0.075 0.068 0.093 0.140   ; 
RECT 0.075 0.140 0.093 0.154   ; 
RECT 0.075 0.154 0.093 0.216   ; 
RECT 0.075 0.216 0.093 0.276   ; 
RECT 0.075 0.276 0.093 0.292   ; 
RECT 0.093 0.140 0.161 0.154   ; 
RECT 0.093 0.276 0.161 0.292   ; 
RECT 0.161 0.140 0.162 0.154   ; 
RECT 0.161 0.154 0.162 0.216   ; 
RECT 0.161 0.276 0.162 0.292   ; 
RECT 0.162 0.140 0.180 0.154   ; 
RECT 0.162 0.154 0.180 0.216   ; 
      LAYER M1 ;
RECT 0.161 0.319 0.351 0.333   ; 
RECT 0.075 0.068 0.093 0.140   ; 
RECT 0.075 0.140 0.093 0.154   ; 
RECT 0.075 0.154 0.093 0.216   ; 
RECT 0.075 0.216 0.093 0.276   ; 
RECT 0.075 0.276 0.093 0.292   ; 
RECT 0.093 0.140 0.161 0.154   ; 
RECT 0.093 0.276 0.161 0.292   ; 
RECT 0.161 0.140 0.162 0.154   ; 
RECT 0.161 0.154 0.162 0.216   ; 
RECT 0.161 0.276 0.162 0.292   ; 
RECT 0.162 0.140 0.180 0.154   ; 
RECT 0.162 0.154 0.180 0.216   ; 
  END
END XOR2_X1

END LIBRARY
#
# End of file
#
