# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2014, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *       NGLibraryCreator, Development_version_64 - build 201405300513        *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on us19.nangate.us for user Lucio Rech (lre).
# Local time is now Tue, 3 Jun 2014, 13:07:07.
# Main process id is 12480.

VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

SITE CORE_TypTyp_0p4_25
  SYMMETRY y ;
  CLASS core ;
  SIZE 0.042 BY 0.504 ;
END CORE_TypTyp_0p4_25



MACRO AND2_X1
  CLASS core ;
  FOREIGN AND2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.252 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.168 0.135187 0.456685 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.0833435 0.0511875 0.34453 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.200812 0.0748125 0.219187 0.42 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.177187 0.522375 ;
  RECT 0.177187 0.485625 0.258562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.258562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0748125 0.106312 0.093122 0.124687 ;
  RECT 0.0748125 0.124687 0.093122 0.280875 ;
  RECT 0.0748125 0.280875 0.093122 0.357 ;
  RECT 0.093122 0.106312 0.158812 0.124687 ;
  RECT 0.158812 0.106312 0.177187 0.124687 ;
  RECT 0.158812 0.124687 0.177187 0.280875 ;
      LAYER M1 ;
  RECT 0.0748125 0.106312 0.093122 0.124687 ;
  RECT 0.0748125 0.124687 0.093122 0.280875 ;
  RECT 0.0748125 0.280875 0.093122 0.357 ;
  RECT 0.093122 0.106312 0.158812 0.124687 ;
  RECT 0.158812 0.106312 0.177187 0.124687 ;
  RECT 0.158812 0.124687 0.177187 0.280875 ;
  END
END AND2_X1

MACRO AND2_X2
  CLASS core ;
  FOREIGN AND2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.252 BY 0.504 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.100 0.168 0.116 0.336   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.025 0.163 0.047 0.341   ; 
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.170 0.042 0.172 0.085   ; 
RECT 0.170 0.419 0.172 0.462   ; 
RECT 0.172 0.042 0.188 0.085   ; 
RECT 0.172 0.085 0.188 0.419   ; 
RECT 0.172 0.419 0.188 0.462   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.006 0.486 0.152 0.522   ; 
RECT 0.152 0.486 0.258 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.006 -0.018 0.258 0.018   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.030 0.377 0.046 0.395   ; 
RECT 0.046 0.109 0.136 0.127   ; 
RECT 0.046 0.377 0.136 0.395   ; 
RECT 0.136 0.109 0.152 0.127   ; 
RECT 0.136 0.127 0.152 0.377   ; 
RECT 0.136 0.377 0.152 0.395   ; 
      LAYER M1 ;
RECT 0.030 0.377 0.046 0.395   ; 
RECT 0.046 0.109 0.136 0.127   ; 
RECT 0.046 0.377 0.136 0.395   ; 
RECT 0.136 0.109 0.152 0.127   ; 
RECT 0.136 0.127 0.152 0.377   ; 
RECT 0.136 0.377 0.152 0.395   ; 
  END
END AND2_X2


MACRO AND3_X1
  CLASS core ;
  FOREIGN AND3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.336 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.200812 0.126 0.219187 0.378 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.113466 0.126 0.138469 0.378 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0315 0.126 0.0525 0.378 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.284813 0.0748125 0.303187 0.429187 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.261188 0.522375 ;
  RECT 0.261188 0.485625 0.342562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.342562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.051844 0.065625 0.156187 0.086625 ;
  RECT 0.0354375 0.414095 0.179812 0.43247 ;
  RECT 0.179812 0.062344 0.242812 0.089906 ;
  RECT 0.179812 0.414095 0.242812 0.43247 ;
  RECT 0.242812 0.062344 0.261188 0.089906 ;
  RECT 0.242812 0.089906 0.261188 0.414095 ;
  RECT 0.242812 0.414095 0.261188 0.43247 ;
      LAYER M1 ;
  RECT 0.051844 0.065625 0.156187 0.086625 ;
  RECT 0.0354375 0.414095 0.179812 0.43247 ;
  RECT 0.179812 0.062344 0.242812 0.089906 ;
  RECT 0.179812 0.414095 0.242812 0.43247 ;
  RECT 0.242812 0.062344 0.261188 0.089906 ;
  RECT 0.242812 0.089906 0.261188 0.414095 ;
  RECT 0.242812 0.414095 0.261188 0.43247 ;
  END
END AND3_X1

MACRO AND3_X2
  CLASS core ;
  FOREIGN AND3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.336 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.21 0.135187 0.336655 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0295312 0.168 0.054469 0.336 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.198187 0.177187 0.352405 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.240187 0.042 0.242812 0.103031 ;
  RECT 0.240187 0.418687 0.242812 0.462 ;
  RECT 0.242812 0.042 0.261188 0.103031 ;
  RECT 0.242812 0.103031 0.261188 0.418687 ;
  RECT 0.242812 0.418687 0.261188 0.462 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.219187 0.522375 ;
  RECT 0.219187 0.485625 0.342562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.342562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0315 0.04725 0.0525 0.102375 ;
  RECT 0.0315 0.102375 0.0525 0.123375 ;
  RECT 0.0525 0.102375 0.195562 0.123375 ;
  RECT 0.0354375 0.38128 0.0958125 0.40228 ;
  RECT 0.0958125 0.147 0.200812 0.165375 ;
  RECT 0.0958125 0.38128 0.200812 0.40228 ;
  RECT 0.200812 0.147 0.219187 0.165375 ;
  RECT 0.200812 0.165375 0.219187 0.38128 ;
  RECT 0.200812 0.38128 0.219187 0.40228 ;
      LAYER M1 ;
  RECT 0.0315 0.04725 0.0525 0.102375 ;
  RECT 0.0315 0.102375 0.0525 0.123375 ;
  RECT 0.0525 0.102375 0.195562 0.123375 ;
  RECT 0.0354375 0.38128 0.0958125 0.40228 ;
  RECT 0.0958125 0.147 0.200812 0.165375 ;
  RECT 0.0958125 0.38128 0.200812 0.40228 ;
  RECT 0.200812 0.147 0.219187 0.165375 ;
  RECT 0.200812 0.165375 0.219187 0.38128 ;
  RECT 0.200812 0.38128 0.219187 0.40228 ;
  END
END AND3_X2

MACRO AND4_X1
  CLASS core ;
  FOREIGN AND4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.378 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.242812 0.126 0.261188 0.378 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.1575 0.126 0.1785 0.378 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.126 0.093122 0.336 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.126 0.0511875 0.378 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.326813 0.0748125 0.345187 0.429187 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.303187 0.522375 ;
  RECT 0.303187 0.485625 0.384562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.384562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0538125 0.417375 0.221812 0.438375 ;
  RECT 0.221812 0.065625 0.284813 0.086625 ;
  RECT 0.221812 0.417375 0.284813 0.438375 ;
  RECT 0.284813 0.065625 0.303187 0.086625 ;
  RECT 0.284813 0.086625 0.303187 0.417375 ;
  RECT 0.284813 0.417375 0.303187 0.438375 ;
  RECT 0.0924655 0.064969 0.195562 0.096469 ;
      LAYER M1 ;
  RECT 0.0538125 0.417375 0.221812 0.438375 ;
  RECT 0.221812 0.065625 0.284813 0.086625 ;
  RECT 0.221812 0.417375 0.284813 0.438375 ;
  RECT 0.284813 0.065625 0.303187 0.086625 ;
  RECT 0.284813 0.086625 0.303187 0.417375 ;
  RECT 0.284813 0.417375 0.303187 0.438375 ;
  RECT 0.0924655 0.064969 0.195562 0.096469 ;
  END
END AND4_X1

MACRO AND4_X2
  CLASS core ;
  FOREIGN AND4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.378 BY 0.504 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
 RECT 0.219 0.158 0.235 0.378   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
 RECT 0.143 0.126 0.159 0.379   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
 RECT 0.067 0.126 0.084 0.379   ; 
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
 RECT 0.030 0.126 0.046 0.379   ; 
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
 RECT 0.294 0.063 0.311 0.420   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
 RECT -0.006 0.486 0.273 0.522   ; 
 RECT 0.273 0.486 0.384 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
 RECT -0.006 -0.018 0.384 0.018   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
 RECT 0.084 0.066 0.176 0.087   ; 
 RECT 0.048 0.417 0.202 0.438   ; 
 RECT 0.202 0.108 0.256 0.129   ; 
 RECT 0.202 0.417 0.256 0.438   ; 
 RECT 0.256 0.108 0.273 0.129   ; 
 RECT 0.256 0.129 0.273 0.417   ; 
 RECT 0.256 0.417 0.273 0.438   ; 
      LAYER M1 ;
 RECT 0.084 0.066 0.176 0.087   ; 
 RECT 0.048 0.417 0.202 0.438   ; 
 RECT 0.202 0.108 0.256 0.129   ; 
 RECT 0.202 0.417 0.256 0.438   ; 
 RECT 0.256 0.108 0.273 0.129   ; 
 RECT 0.256 0.129 0.273 0.417   ; 
 RECT 0.256 0.417 0.273 0.438   ; 
  END
END AND4_X2

MACRO ANTENNA
  CLASS core ;
  FOREIGN ANTENNA 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.126 BY 0.504 ;
END ANTENNA

MACRO AOI21_X1
  CLASS core ;
  FOREIGN AOI21_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.252 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.126 0.135187 0.336 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.0879375 0.0511875 0.336 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.200812 0.126 0.219187 0.336 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.065625 0.093122 0.086625 ;
  RECT 0.0748125 0.086625 0.093122 0.35175 ;
  RECT 0.093122 0.065625 0.200812 0.086625 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.195562 0.522375 ;
  RECT 0.195562 0.485625 0.258562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.258562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0315 0.380625 0.0525 0.401625 ;
  RECT 0.0315 0.401625 0.0525 0.462 ;
  RECT 0.0525 0.380625 0.195562 0.401625 ;
      LAYER M1 ;
  RECT 0.0315 0.380625 0.0525 0.401625 ;
  RECT 0.0315 0.401625 0.0525 0.462 ;
  RECT 0.0525 0.380625 0.195562 0.401625 ;
  END
END AOI21_X1

MACRO AOI21_X2
  CLASS core ;
  FOREIGN AOI21_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
 SIZE 0.252 BY 0.504 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
 RECT 0.162 0.198 0.174 0.294   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
 RECT 0.106 0.151 0.118 0.169   ; 
 RECT 0.106 0.169 0.118 0.294   ; 
 RECT 0.106 0.294 0.118 0.336   ; 
 RECT 0.118 0.151 0.216 0.169   ; 
 RECT 0.216 0.151 0.232 0.169   ; 
 RECT 0.216 0.169 0.232 0.294   ; 
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
 RECT 0.050 0.168 0.062 0.294   ; 
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
 RECT 0.034 0.109 0.078 0.127   ; 
 RECT 0.078 0.109 0.090 0.127   ; 
 RECT 0.078 0.127 0.090 0.321   ; 
 RECT 0.078 0.321 0.090 0.375   ; 
 RECT 0.078 0.375 0.090 0.393   ; 
 RECT 0.090 0.109 0.188 0.127   ; 
 RECT 0.090 0.375 0.188 0.393   ; 
 RECT 0.188 0.375 0.190 0.393   ; 
 RECT 0.190 0.321 0.202 0.375   ; 
 RECT 0.190 0.375 0.202 0.393   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
 RECT -0.004 0.486 0.230 0.522   ; 
 RECT 0.230 0.486 0.234 0.522   ; 
 RECT 0.234 0.486 0.256 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
 RECT -0.004 -0.018 0.256 0.018   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
 RECT 0.021 0.361 0.035 0.417   ; 
 RECT 0.021 0.417 0.035 0.439   ; 
 RECT 0.035 0.417 0.218 0.439   ; 
 RECT 0.218 0.339 0.230 0.361   ; 
 RECT 0.218 0.361 0.230 0.417   ; 
 RECT 0.218 0.417 0.230 0.439   ; 
 RECT 0.064 0.067 0.234 0.085   ; 
      LAYER M1 ;
 RECT 0.021 0.361 0.035 0.417   ; 
 RECT 0.021 0.417 0.035 0.439   ; 
 RECT 0.035 0.417 0.218 0.439   ; 
 RECT 0.218 0.339 0.230 0.361   ; 
 RECT 0.218 0.361 0.230 0.417   ; 
 RECT 0.218 0.417 0.230 0.439   ; 
 RECT 0.064 0.067 0.234 0.085   ; 
  END
END AOI21_X2

MACRO AOI22_X1
  CLASS core ;
  FOREIGN AOI22_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.294 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.126 0.177187 0.336 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.242812 0.126 0.261188 0.31828 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.129937 0.093122 0.378 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.126 0.0511875 0.378 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0924655 0.066872 0.200812 0.0853125 ;
  RECT 0.200812 0.066872 0.219187 0.0853125 ;
  RECT 0.200812 0.0853125 0.219187 0.381937 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.261188 0.522375 ;
  RECT 0.261188 0.485625 0.300563 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.300563 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0538125 0.413438 0.242812 0.442312 ;
  RECT 0.242812 0.362905 0.261188 0.413438 ;
  RECT 0.242812 0.413438 0.261188 0.442312 ;
      LAYER M1 ;
  RECT 0.0538125 0.413438 0.242812 0.442312 ;
  RECT 0.242812 0.362905 0.261188 0.413438 ;
  RECT 0.242812 0.413438 0.261188 0.442312 ;
  END
END AOI22_X1

MACRO AOI22_X2
  CLASS core ;
  FOREIGN AOI22_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
 SIZE 0.294 BY 0.504 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
 RECT 0.166 0.180 0.177 0.198   ; 
 RECT 0.166 0.198 0.177 0.321   ; 
 RECT 0.166 0.321 0.177 0.336   ; 
 RECT 0.177 0.180 0.250 0.198   ; 
 RECT 0.250 0.180 0.264 0.198   ; 
 RECT 0.264 0.180 0.275 0.198   ; 
 RECT 0.264 0.198 0.275 0.321   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
 RECT 0.215 0.243 0.226 0.336   ; 
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
 RECT 0.117 0.201 0.128 0.345   ; 
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
 RECT 0.019 0.159 0.030 0.336   ; 
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
 RECT 0.093 0.131 0.103 0.150   ; 
 RECT 0.093 0.150 0.103 0.150   ; 
 RECT 0.093 0.150 0.103 0.210   ; 
 RECT 0.103 0.131 0.139 0.150   ; 
 RECT 0.139 0.131 0.142 0.150   ; 
 RECT 0.142 0.131 0.152 0.150   ; 
 RECT 0.142 0.150 0.152 0.150   ; 
 RECT 0.142 0.150 0.152 0.210   ; 
 RECT 0.142 0.210 0.152 0.304   ; 
 RECT 0.142 0.304 0.152 0.373   ; 
 RECT 0.142 0.373 0.152 0.395   ; 
 RECT 0.152 0.131 0.240 0.150   ; 
 RECT 0.152 0.150 0.240 0.150   ; 
 RECT 0.152 0.373 0.240 0.395   ; 
 RECT 0.240 0.131 0.250 0.150   ; 
 RECT 0.240 0.150 0.250 0.150   ; 
 RECT 0.240 0.304 0.250 0.373   ; 
 RECT 0.240 0.373 0.250 0.395   ; 
 RECT 0.250 0.131 0.264 0.150   ; 
 RECT 0.250 0.150 0.264 0.150   ; 
 RECT 0.264 0.063 0.275 0.131   ; 
 RECT 0.264 0.131 0.275 0.150   ; 
 RECT 0.264 0.150 0.275 0.150   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
 RECT -0.004 0.486 0.275 0.522   ; 
 RECT 0.275 0.486 0.298 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
 RECT -0.004 -0.018 0.298 0.018   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
 RECT 0.155 0.087 0.240 0.108   ; 
 RECT 0.240 0.047 0.250 0.087   ; 
 RECT 0.240 0.087 0.250 0.108   ; 
 RECT 0.029 0.419 0.264 0.437   ; 
 RECT 0.264 0.366 0.275 0.419   ; 
 RECT 0.264 0.419 0.275 0.437   ; 
 RECT 0.033 0.057 0.139 0.095   ; 
      LAYER M1 ;
 RECT 0.155 0.087 0.240 0.108   ; 
 RECT 0.240 0.047 0.250 0.087   ; 
 RECT 0.240 0.087 0.250 0.108   ; 
 RECT 0.029 0.419 0.264 0.437   ; 
 RECT 0.264 0.366 0.275 0.419   ; 
 RECT 0.264 0.419 0.275 0.437   ; 
 RECT 0.033 0.057 0.139 0.095   ; 
  END
END AOI22_X2

MACRO BUF_X1
  CLASS core ;
  FOREIGN BUF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.21 BY 0.504 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.126 0.0511875 0.378 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.1575 0.0748125 0.1785 0.462 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.093778 0.522375 ;
  RECT 0.093778 0.485625 0.216562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.216562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0748125 0.04725 0.075469 0.121406 ;
  RECT 0.0748125 0.121406 0.075469 0.139781 ;
  RECT 0.0748125 0.280875 0.075469 0.29925 ;
  RECT 0.0748125 0.29925 0.075469 0.366187 ;
  RECT 0.075469 0.04725 0.093122 0.121406 ;
  RECT 0.075469 0.121406 0.093122 0.139781 ;
  RECT 0.075469 0.139781 0.093122 0.280875 ;
  RECT 0.075469 0.280875 0.093122 0.29925 ;
  RECT 0.075469 0.29925 0.093122 0.366187 ;
  RECT 0.093122 0.121406 0.093778 0.139781 ;
  RECT 0.093122 0.139781 0.093778 0.280875 ;
  RECT 0.093122 0.280875 0.093778 0.29925 ;
      LAYER M1 ;
  RECT 0.0748125 0.04725 0.075469 0.121406 ;
  RECT 0.0748125 0.121406 0.075469 0.139781 ;
  RECT 0.0748125 0.280875 0.075469 0.29925 ;
  RECT 0.0748125 0.29925 0.075469 0.366187 ;
  RECT 0.075469 0.04725 0.093122 0.121406 ;
  RECT 0.075469 0.121406 0.093122 0.139781 ;
  RECT 0.075469 0.139781 0.093122 0.280875 ;
  RECT 0.075469 0.280875 0.093122 0.29925 ;
  RECT 0.075469 0.29925 0.093122 0.366187 ;
  RECT 0.093122 0.121406 0.093778 0.139781 ;
  RECT 0.093122 0.139781 0.093778 0.280875 ;
  RECT 0.093122 0.280875 0.093778 0.29925 ;
  END
END BUF_X1

MACRO BUF_X2
  CLASS core ;
  FOREIGN BUF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.21 BY 0.504 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.175219 0.0511875 0.336 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.114122 0.39572 0.116156 0.462 ;
  RECT 0.116156 0.04725 0.116812 0.086625 ;
  RECT 0.116156 0.39572 0.116812 0.462 ;
  RECT 0.116812 0.04725 0.135187 0.086625 ;
  RECT 0.116812 0.086625 0.135187 0.39572 ;
  RECT 0.116812 0.39572 0.135187 0.462 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.093122 0.522375 ;
  RECT 0.093122 0.485625 0.216562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.216562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0275625 0.364875 0.0328125 0.38325 ;
  RECT 0.0275625 0.38325 0.0328125 0.450188 ;
  RECT 0.0328125 0.063 0.0511875 0.126 ;
  RECT 0.0328125 0.126 0.0511875 0.144375 ;
  RECT 0.0328125 0.364875 0.0511875 0.38325 ;
  RECT 0.0328125 0.38325 0.0511875 0.450188 ;
  RECT 0.0511875 0.126 0.056372 0.144375 ;
  RECT 0.0511875 0.364875 0.056372 0.38325 ;
  RECT 0.0511875 0.38325 0.056372 0.450188 ;
  RECT 0.056372 0.126 0.0748125 0.144375 ;
  RECT 0.056372 0.364875 0.0748125 0.38325 ;
  RECT 0.0748125 0.126 0.093122 0.144375 ;
  RECT 0.0748125 0.144375 0.093122 0.364875 ;
  RECT 0.0748125 0.364875 0.093122 0.38325 ;
      LAYER M1 ;
  RECT 0.0275625 0.364875 0.0328125 0.38325 ;
  RECT 0.0275625 0.38325 0.0328125 0.450188 ;
  RECT 0.0328125 0.063 0.0511875 0.126 ;
  RECT 0.0328125 0.126 0.0511875 0.144375 ;
  RECT 0.0328125 0.364875 0.0511875 0.38325 ;
  RECT 0.0328125 0.38325 0.0511875 0.450188 ;
  RECT 0.0511875 0.126 0.056372 0.144375 ;
  RECT 0.0511875 0.364875 0.056372 0.38325 ;
  RECT 0.0511875 0.38325 0.056372 0.450188 ;
  RECT 0.056372 0.126 0.0748125 0.144375 ;
  RECT 0.056372 0.364875 0.0748125 0.38325 ;
  RECT 0.0748125 0.126 0.093122 0.144375 ;
  RECT 0.0748125 0.144375 0.093122 0.364875 ;
  RECT 0.0748125 0.364875 0.093122 0.38325 ;
  END
END BUF_X2

MACRO BUF_X4
  CLASS core ;
  FOREIGN BUF_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
 SIZE 0.210 BY 0.504 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
 RECT 0.073 0.159 0.084 0.345   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
 RECT 0.059 0.067 0.086 0.085   ; 
 RECT 0.086 0.067 0.111 0.085   ; 
 RECT 0.086 0.419 0.111 0.437   ; 
 RECT 0.111 0.067 0.151 0.085   ; 
 RECT 0.111 0.419 0.151 0.437   ; 
 RECT 0.151 0.067 0.164 0.085   ; 
 RECT 0.151 0.085 0.164 0.419   ; 
 RECT 0.151 0.419 0.164 0.437   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
 RECT -0.004 0.486 0.111 0.522   ; 
 RECT 0.111 0.486 0.214 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
 RECT -0.004 -0.018 0.214 0.018   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
 RECT 0.011 0.109 0.035 0.130   ; 
 RECT 0.035 0.109 0.099 0.130   ; 
 RECT 0.035 0.374 0.099 0.395   ; 
 RECT 0.099 0.109 0.111 0.130   ; 
 RECT 0.099 0.130 0.111 0.374   ; 
 RECT 0.099 0.374 0.111 0.395   ; 
      LAYER M1 ;
 RECT 0.011 0.109 0.035 0.130   ; 
 RECT 0.035 0.109 0.099 0.130   ; 
 RECT 0.035 0.374 0.099 0.395   ; 
 RECT 0.099 0.109 0.111 0.130   ; 
 RECT 0.099 0.130 0.111 0.374   ; 
 RECT 0.099 0.374 0.111 0.395   ; 
  END
END BUF_X4

MACRO BUF_X8
  CLASS core ;
  FOREIGN BUF_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
 SIZE 0.210 BY 0.504 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
 RECT 0.012 0.168 0.018 0.240   ; 
 RECT 0.012 0.240 0.018 0.261   ; 
 RECT 0.012 0.261 0.018 0.336   ; 
 RECT 0.018 0.240 0.070 0.261   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
 RECT 0.079 0.067 0.164 0.085   ; 
 RECT 0.079 0.419 0.164 0.437   ; 
 RECT 0.164 0.067 0.177 0.085   ; 
 RECT 0.164 0.419 0.177 0.437   ; 
 RECT 0.177 0.067 0.183 0.085   ; 
 RECT 0.177 0.085 0.183 0.419   ; 
 RECT 0.177 0.419 0.183 0.437   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
 RECT -0.002 0.486 0.164 0.522   ; 
 RECT 0.164 0.486 0.212 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
 RECT -0.002 -0.018 0.212 0.018   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
 RECT 0.023 0.064 0.027 0.122   ; 
 RECT 0.023 0.122 0.027 0.140   ; 
 RECT 0.027 0.064 0.033 0.122   ; 
 RECT 0.027 0.122 0.033 0.140   ; 
 RECT 0.027 0.346 0.033 0.383   ; 
 RECT 0.027 0.383 0.033 0.440   ; 
 RECT 0.033 0.064 0.037 0.122   ; 
 RECT 0.033 0.122 0.037 0.140   ; 
 RECT 0.033 0.346 0.037 0.383   ; 
 RECT 0.037 0.122 0.083 0.140   ; 
 RECT 0.037 0.346 0.083 0.383   ; 
 RECT 0.083 0.122 0.090 0.140   ; 
 RECT 0.083 0.140 0.090 0.224   ; 
 RECT 0.083 0.224 0.090 0.242   ; 
 RECT 0.083 0.242 0.090 0.346   ; 
 RECT 0.083 0.346 0.090 0.383   ; 
 RECT 0.090 0.224 0.164 0.242   ; 
      LAYER M1 ;
 RECT 0.023 0.064 0.027 0.122   ; 
 RECT 0.023 0.122 0.027 0.140   ; 
 RECT 0.027 0.064 0.033 0.122   ; 
 RECT 0.027 0.122 0.033 0.140   ; 
 RECT 0.027 0.346 0.033 0.383   ; 
 RECT 0.027 0.383 0.033 0.440   ; 
 RECT 0.033 0.064 0.037 0.122   ; 
 RECT 0.033 0.122 0.037 0.140   ; 
 RECT 0.033 0.346 0.037 0.383   ; 
 RECT 0.037 0.122 0.083 0.140   ; 
 RECT 0.037 0.346 0.083 0.383   ; 
 RECT 0.083 0.122 0.090 0.140   ; 
 RECT 0.083 0.140 0.090 0.224   ; 
 RECT 0.083 0.224 0.090 0.242   ; 
 RECT 0.083 0.242 0.090 0.346   ; 
 RECT 0.083 0.346 0.090 0.383   ; 
 RECT 0.090 0.224 0.164 0.242   ; 
  END
END BUF_X8

MACRO BUF_X12
  CLASS core ;
  FOREIGN BUF_X12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
 SIZE 0.294 BY 0.504 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
 RECT 0.010 0.155 0.017 0.240   ; 
 RECT 0.010 0.240 0.017 0.261   ; 
 RECT 0.010 0.261 0.017 0.338   ; 
 RECT 0.017 0.240 0.093 0.261   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
 RECT 0.102 0.067 0.234 0.085   ; 
 RECT 0.102 0.419 0.234 0.437   ; 
 RECT 0.234 0.067 0.248 0.085   ; 
 RECT 0.234 0.419 0.248 0.437   ; 
 RECT 0.248 0.067 0.255 0.085   ; 
 RECT 0.248 0.085 0.255 0.419   ; 
 RECT 0.248 0.419 0.255 0.437   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
 RECT -0.002 0.486 0.234 0.522   ; 
 RECT 0.234 0.486 0.282 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
 RECT -0.002 -0.018 0.282 0.018   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
 RECT 0.021 0.362 0.024 0.383   ; 
 RECT 0.021 0.383 0.024 0.440   ; 
 RECT 0.024 0.064 0.031 0.121   ; 
 RECT 0.024 0.121 0.031 0.142   ; 
 RECT 0.024 0.362 0.031 0.383   ; 
 RECT 0.024 0.383 0.031 0.440   ; 
 RECT 0.031 0.121 0.034 0.142   ; 
 RECT 0.031 0.362 0.034 0.383   ; 
 RECT 0.031 0.383 0.034 0.440   ; 
 RECT 0.034 0.121 0.101 0.142   ; 
 RECT 0.034 0.362 0.101 0.383   ; 
 RECT 0.101 0.121 0.107 0.142   ; 
 RECT 0.101 0.142 0.107 0.243   ; 
 RECT 0.101 0.243 0.107 0.261   ; 
 RECT 0.101 0.261 0.107 0.362   ; 
 RECT 0.101 0.362 0.107 0.383   ; 
 RECT 0.107 0.243 0.234 0.261   ; 
      LAYER M1 ;
 RECT 0.021 0.362 0.024 0.383   ; 
 RECT 0.021 0.383 0.024 0.440   ; 
 RECT 0.024 0.064 0.031 0.121   ; 
 RECT 0.024 0.121 0.031 0.142   ; 
 RECT 0.024 0.362 0.031 0.383   ; 
 RECT 0.024 0.383 0.031 0.440   ; 
 RECT 0.031 0.121 0.034 0.142   ; 
 RECT 0.031 0.362 0.034 0.383   ; 
 RECT 0.031 0.383 0.034 0.440   ; 
 RECT 0.034 0.121 0.101 0.142   ; 
 RECT 0.034 0.362 0.101 0.383   ; 
 RECT 0.101 0.121 0.107 0.142   ; 
 RECT 0.101 0.142 0.107 0.243   ; 
 RECT 0.101 0.243 0.107 0.261   ; 
 RECT 0.101 0.261 0.107 0.362   ; 
 RECT 0.101 0.362 0.107 0.383   ; 
 RECT 0.107 0.243 0.234 0.261   ; 
  END
END BUF_X12


MACRO BUF_X16
  CLASS core ;
  FOREIGN BUF_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
 SIZE 0.294 BY 0.504 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
 RECT 0.008 0.152 0.013 0.233   ; 
 RECT 0.008 0.233 0.013 0.271   ; 
 RECT 0.008 0.271 0.013 0.336   ; 
 RECT 0.013 0.233 0.093 0.271   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
 RECT 0.100 0.067 0.245 0.085   ; 
 RECT 0.100 0.415 0.245 0.433   ; 
 RECT 0.245 0.067 0.256 0.085   ; 
 RECT 0.245 0.415 0.256 0.433   ; 
 RECT 0.256 0.067 0.261 0.085   ; 
 RECT 0.256 0.085 0.261 0.415   ; 
 RECT 0.256 0.415 0.261 0.433   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
 RECT -0.002 0.486 0.245 0.522   ; 
 RECT 0.245 0.486 0.282 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
 RECT -0.002 -0.018 0.282 0.018   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
 RECT 0.019 0.064 0.024 0.135   ; 
 RECT 0.019 0.135 0.024 0.153   ; 
 RECT 0.019 0.301 0.024 0.319   ; 
 RECT 0.019 0.319 0.024 0.422   ; 
 RECT 0.024 0.135 0.099 0.153   ; 
 RECT 0.024 0.301 0.099 0.319   ; 
 RECT 0.099 0.135 0.104 0.153   ; 
 RECT 0.099 0.153 0.104 0.241   ; 
 RECT 0.099 0.241 0.104 0.260   ; 
 RECT 0.099 0.260 0.104 0.301   ; 
 RECT 0.099 0.301 0.104 0.319   ; 
 RECT 0.104 0.241 0.245 0.260   ; 
      LAYER M1 ;
 RECT 0.019 0.064 0.024 0.135   ; 
 RECT 0.019 0.135 0.024 0.153   ; 
 RECT 0.019 0.301 0.024 0.319   ; 
 RECT 0.019 0.319 0.024 0.422   ; 
 RECT 0.024 0.135 0.099 0.153   ; 
 RECT 0.024 0.301 0.099 0.319   ; 
 RECT 0.099 0.135 0.104 0.153   ; 
 RECT 0.099 0.153 0.104 0.241   ; 
 RECT 0.099 0.241 0.104 0.260   ; 
 RECT 0.099 0.260 0.104 0.301   ; 
 RECT 0.099 0.301 0.104 0.319   ; 
 RECT 0.104 0.241 0.245 0.260   ; 
  END
END BUF_X16

MACRO CLKBUF_X1
  CLASS core ;
  FOREIGN CLKBUF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.21 BY 0.504 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.126 0.0511875 0.378 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.1575 0.0748125 0.1785 0.462 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.093778 0.522375 ;
  RECT 0.093778 0.485625 0.216562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.216562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0748125 0.04725 0.075469 0.121406 ;
  RECT 0.0748125 0.121406 0.075469 0.139781 ;
  RECT 0.0748125 0.257905 0.075469 0.300563 ;
  RECT 0.0748125 0.300563 0.075469 0.34322 ;
  RECT 0.075469 0.04725 0.093122 0.121406 ;
  RECT 0.075469 0.121406 0.093122 0.139781 ;
  RECT 0.075469 0.139781 0.093122 0.257905 ;
  RECT 0.075469 0.257905 0.093122 0.300563 ;
  RECT 0.075469 0.300563 0.093122 0.34322 ;
  RECT 0.093122 0.121406 0.093778 0.139781 ;
  RECT 0.093122 0.139781 0.093778 0.257905 ;
  RECT 0.093122 0.257905 0.093778 0.300563 ;
      LAYER M1 ;
  RECT 0.0748125 0.04725 0.075469 0.121406 ;
  RECT 0.0748125 0.121406 0.075469 0.139781 ;
  RECT 0.0748125 0.257905 0.075469 0.300563 ;
  RECT 0.0748125 0.300563 0.075469 0.34322 ;
  RECT 0.075469 0.04725 0.093122 0.121406 ;
  RECT 0.075469 0.121406 0.093122 0.139781 ;
  RECT 0.075469 0.139781 0.093122 0.257905 ;
  RECT 0.075469 0.257905 0.093122 0.300563 ;
  RECT 0.075469 0.300563 0.093122 0.34322 ;
  RECT 0.093122 0.121406 0.093778 0.139781 ;
  RECT 0.093122 0.139781 0.093778 0.257905 ;
  RECT 0.093122 0.257905 0.093778 0.300563 ;
  END
END CLKBUF_X1

MACRO CLKBUF_X2
  CLASS core ;
  FOREIGN CLKBUF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.21 BY 0.504 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.19425 0.0511875 0.336 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.114122 0.418687 0.116812 0.462 ;
  RECT 0.116812 0.04725 0.135187 0.418687 ;
  RECT 0.116812 0.418687 0.135187 0.462 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.093122 0.522375 ;
  RECT 0.093122 0.485625 0.216562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.216562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0315 0.0846565 0.0525 0.126 ;
  RECT 0.0315 0.126 0.0525 0.144375 ;
  RECT 0.0315 0.364875 0.0525 0.38325 ;
  RECT 0.0315 0.38325 0.0525 0.450188 ;
  RECT 0.0525 0.126 0.0748125 0.144375 ;
  RECT 0.0525 0.364875 0.0748125 0.38325 ;
  RECT 0.0748125 0.126 0.093122 0.144375 ;
  RECT 0.0748125 0.144375 0.093122 0.364875 ;
  RECT 0.0748125 0.364875 0.093122 0.38325 ;
      LAYER M1 ;
  RECT 0.0315 0.0846565 0.0525 0.126 ;
  RECT 0.0315 0.126 0.0525 0.144375 ;
  RECT 0.0315 0.364875 0.0525 0.38325 ;
  RECT 0.0315 0.38325 0.0525 0.450188 ;
  RECT 0.0525 0.126 0.0748125 0.144375 ;
  RECT 0.0525 0.364875 0.0748125 0.38325 ;
  RECT 0.0748125 0.126 0.093122 0.144375 ;
  RECT 0.0748125 0.144375 0.093122 0.364875 ;
  RECT 0.0748125 0.364875 0.093122 0.38325 ;
  END
END CLKBUF_X2

MACRO CLKBUF_X4
  CLASS core ;
  FOREIGN CLKBUF_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
 SIZE 0.210 BY 0.504 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
 RECT 0.047 0.159 0.058 0.345   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
 RECT 0.059 0.067 0.084 0.085   ; 
 RECT 0.084 0.067 0.084 0.085   ; 
 RECT 0.084 0.419 0.084 0.437   ; 
 RECT 0.084 0.067 0.151 0.085   ; 
 RECT 0.084 0.419 0.151 0.437   ; 
 RECT 0.151 0.067 0.164 0.085   ; 
 RECT 0.151 0.085 0.164 0.419   ; 
 RECT 0.151 0.419 0.164 0.437   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
 RECT -0.004 0.486 0.084 0.522   ; 
 RECT 0.084 0.486 0.214 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
 RECT -0.004 -0.018 0.214 0.018   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
 RECT 0.017 0.109 0.034 0.127   ; 
 RECT 0.034 0.109 0.073 0.127   ; 
 RECT 0.034 0.377 0.073 0.395   ; 
 RECT 0.073 0.109 0.084 0.127   ; 
 RECT 0.073 0.127 0.084 0.377   ; 
 RECT 0.073 0.377 0.084 0.395   ; 
      LAYER M1 ;
 RECT 0.017 0.109 0.034 0.127   ; 
 RECT 0.034 0.109 0.073 0.127   ; 
 RECT 0.034 0.377 0.073 0.395   ; 
 RECT 0.073 0.109 0.084 0.127   ; 
 RECT 0.073 0.127 0.084 0.377   ; 
 RECT 0.073 0.377 0.084 0.395   ; 
  END
END CLKBUF_X4

MACRO CLKBUF_X8
  CLASS core ;
  FOREIGN CLKBUF_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
 SIZE 0.210 BY 0.504 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
 RECT 0.012 0.168 0.018 0.215   ; 
 RECT 0.012 0.215 0.018 0.234   ; 
 RECT 0.012 0.234 0.018 0.336   ; 
 RECT 0.018 0.168 0.019 0.215   ; 
 RECT 0.018 0.215 0.019 0.234   ; 
 RECT 0.019 0.215 0.075 0.234   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
 RECT 0.079 0.067 0.168 0.085   ; 
 RECT 0.079 0.419 0.168 0.437   ; 
 RECT 0.168 0.067 0.177 0.085   ; 
 RECT 0.168 0.419 0.177 0.437   ; 
 RECT 0.177 0.067 0.183 0.085   ; 
 RECT 0.177 0.085 0.183 0.419   ; 
 RECT 0.177 0.419 0.183 0.437   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
 RECT -0.002 0.486 0.168 0.522   ; 
 RECT 0.168 0.486 0.212 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
 RECT -0.002 -0.018 0.212 0.018   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
 RECT 0.012 0.109 0.027 0.127   ; 
 RECT 0.027 0.109 0.033 0.127   ; 
 RECT 0.027 0.295 0.033 0.316   ; 
 RECT 0.027 0.316 0.033 0.356   ; 
 RECT 0.033 0.109 0.095 0.127   ; 
 RECT 0.033 0.295 0.095 0.316   ; 
 RECT 0.095 0.109 0.102 0.127   ; 
 RECT 0.095 0.127 0.102 0.234   ; 
 RECT 0.095 0.234 0.102 0.272   ; 
 RECT 0.095 0.272 0.102 0.295   ; 
 RECT 0.095 0.295 0.102 0.316   ; 
 RECT 0.102 0.234 0.168 0.272   ; 
      LAYER M1 ;
 RECT 0.012 0.109 0.027 0.127   ; 
 RECT 0.027 0.109 0.033 0.127   ; 
 RECT 0.027 0.295 0.033 0.316   ; 
 RECT 0.027 0.316 0.033 0.356   ; 
 RECT 0.033 0.109 0.095 0.127   ; 
 RECT 0.033 0.295 0.095 0.316   ; 
 RECT 0.095 0.109 0.102 0.127   ; 
 RECT 0.095 0.127 0.102 0.234   ; 
 RECT 0.095 0.234 0.102 0.272   ; 
 RECT 0.095 0.272 0.102 0.295   ; 
 RECT 0.095 0.295 0.102 0.316   ; 
 RECT 0.102 0.234 0.168 0.272   ; 
  END
END CLKBUF_X8

MACRO CLKBUF_X12
  CLASS core ;
  FOREIGN CLKBUF_X12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
 SIZE 0.294 BY 0.504 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
 RECT 0.010 0.156 0.018 0.221   ; 
 RECT 0.010 0.221 0.018 0.241   ; 
 RECT 0.010 0.241 0.018 0.348   ; 
 RECT 0.018 0.221 0.093 0.241   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
 RECT 0.102 0.067 0.218 0.085   ; 
 RECT 0.102 0.419 0.218 0.437   ; 
 RECT 0.218 0.067 0.248 0.085   ; 
 RECT 0.218 0.419 0.248 0.437   ; 
 RECT 0.248 0.067 0.255 0.085   ; 
 RECT 0.248 0.085 0.255 0.419   ; 
 RECT 0.248 0.419 0.255 0.437   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
 RECT -0.002 0.486 0.218 0.522   ; 
 RECT 0.218 0.486 0.282 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
 RECT -0.002 -0.018 0.282 0.018   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
 RECT 0.009 0.109 0.025 0.127   ; 
 RECT 0.025 0.109 0.031 0.127   ; 
 RECT 0.025 0.361 0.031 0.379   ; 
 RECT 0.025 0.379 0.031 0.440   ; 
 RECT 0.031 0.109 0.101 0.127   ; 
 RECT 0.031 0.361 0.101 0.379   ; 
 RECT 0.101 0.109 0.107 0.127   ; 
 RECT 0.101 0.127 0.107 0.206   ; 
 RECT 0.101 0.206 0.107 0.227   ; 
 RECT 0.101 0.227 0.107 0.361   ; 
 RECT 0.101 0.361 0.107 0.379   ; 
 RECT 0.107 0.109 0.108 0.127   ; 
 RECT 0.107 0.127 0.108 0.206   ; 
 RECT 0.107 0.206 0.108 0.227   ; 
 RECT 0.108 0.206 0.218 0.227   ; 
      LAYER M1 ;
 RECT 0.009 0.109 0.025 0.127   ; 
 RECT 0.025 0.109 0.031 0.127   ; 
 RECT 0.025 0.361 0.031 0.379   ; 
 RECT 0.025 0.379 0.031 0.440   ; 
 RECT 0.031 0.109 0.101 0.127   ; 
 RECT 0.031 0.361 0.101 0.379   ; 
 RECT 0.101 0.109 0.107 0.127   ; 
 RECT 0.101 0.127 0.107 0.206   ; 
 RECT 0.101 0.206 0.107 0.227   ; 
 RECT 0.101 0.227 0.107 0.361   ; 
 RECT 0.101 0.361 0.107 0.379   ; 
 RECT 0.107 0.109 0.108 0.127   ; 
 RECT 0.107 0.127 0.108 0.206   ; 
 RECT 0.107 0.206 0.108 0.227   ; 
 RECT 0.108 0.206 0.218 0.227   ; 
  END
END CLKBUF_X12

MACRO CLKBUF_X16
  CLASS core ;
  FOREIGN CLKBUF_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
 SIZE 0.294 BY 0.504 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
 RECT 0.008 0.146 0.013 0.214   ; 
 RECT 0.008 0.214 0.013 0.235   ; 
 RECT 0.008 0.235 0.013 0.345   ; 
 RECT 0.013 0.214 0.093 0.235   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
 RECT 0.100 0.057 0.245 0.095   ; 
 RECT 0.100 0.409 0.245 0.447   ; 
 RECT 0.245 0.057 0.256 0.095   ; 
 RECT 0.245 0.409 0.256 0.447   ; 
 RECT 0.256 0.057 0.261 0.095   ; 
 RECT 0.256 0.095 0.261 0.409   ; 
 RECT 0.256 0.409 0.261 0.447   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
 RECT -0.002 0.486 0.245 0.522   ; 
 RECT 0.245 0.486 0.282 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
 RECT -0.002 -0.018 0.282 0.018   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
 RECT 0.019 0.072 0.024 0.135   ; 
 RECT 0.019 0.135 0.024 0.153   ; 
 RECT 0.019 0.345 0.024 0.369   ; 
 RECT 0.019 0.369 0.024 0.419   ; 
 RECT 0.024 0.135 0.100 0.153   ; 
 RECT 0.024 0.345 0.100 0.369   ; 
 RECT 0.100 0.135 0.110 0.153   ; 
 RECT 0.100 0.153 0.110 0.207   ; 
 RECT 0.100 0.207 0.110 0.226   ; 
 RECT 0.100 0.226 0.110 0.345   ; 
 RECT 0.100 0.345 0.110 0.369   ; 
 RECT 0.110 0.207 0.245 0.226   ; 
      LAYER M1 ;
 RECT 0.019 0.072 0.024 0.135   ; 
 RECT 0.019 0.135 0.024 0.153   ; 
 RECT 0.019 0.345 0.024 0.369   ; 
 RECT 0.019 0.369 0.024 0.419   ; 
 RECT 0.024 0.135 0.100 0.153   ; 
 RECT 0.024 0.345 0.100 0.369   ; 
 RECT 0.100 0.135 0.110 0.153   ; 
 RECT 0.100 0.153 0.110 0.207   ; 
 RECT 0.100 0.207 0.110 0.226   ; 
 RECT 0.100 0.226 0.110 0.345   ; 
 RECT 0.100 0.345 0.110 0.369   ; 
 RECT 0.110 0.207 0.245 0.226   ; 
  END
END CLKBUF_X16

MACRO DFFRNQ_X1
  CLASS core ;
  FOREIGN DFFRNQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 1.092 BY 0.504 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.158812 0.177187 0.345187 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
  RECT 0.462 0.179812 0.744125 0.198187 ;
  RECT 0.744125 0.179812 0.87019 0.198187 ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.168 0.0511875 0.336 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 1.0395 0.042 1.0605 0.462 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.093122 0.522375 ;
  RECT 0.093122 0.485625 0.135187 0.522375 ;
  RECT 0.135187 0.485625 0.219187 0.522375 ;
  RECT 0.219187 0.485625 0.261188 0.522375 ;
  RECT 0.261188 0.485625 0.345187 0.522375 ;
  RECT 0.345187 0.485625 0.53412 0.522375 ;
  RECT 0.53412 0.485625 0.597185 0.522375 ;
  RECT 0.597185 0.485625 0.63919 0.522375 ;
  RECT 0.63919 0.485625 0.723185 0.522375 ;
  RECT 0.723185 0.485625 0.779625 0.522375 ;
  RECT 0.779625 0.485625 0.9765 0.522375 ;
  RECT 0.9765 0.485625 1.09856 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 1.09856 0.018375 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
  RECT 0.0958125 0.137812 0.744125 0.156187 ;
  RECT 0.0538125 0.347813 0.744125 0.366187 ;
      LAYER MINT1 ;
  RECT 0.0958125 0.137812 0.744125 0.156187 ;
  RECT 0.0538125 0.347813 0.744125 0.366187 ;
      LAYER M1 ;
  RECT 0.116812 0.04725 0.135187 0.456685 ;
  RECT 0.200812 0.04725 0.219187 0.456685 ;
  RECT 0.347813 0.408845 0.53412 0.446905 ;
  RECT 0.284813 0.066872 0.303187 0.0853125 ;
  RECT 0.284813 0.0853125 0.303187 0.287438 ;
  RECT 0.284813 0.287438 0.303187 0.439688 ;
  RECT 0.303187 0.066872 0.525 0.0853125 ;
  RECT 0.525 0.066872 0.543375 0.0853125 ;
  RECT 0.525 0.0853125 0.543375 0.287438 ;
  RECT 0.378 0.216562 0.396375 0.332062 ;
  RECT 0.378 0.332062 0.396375 0.350438 ;
  RECT 0.396375 0.332062 0.57881 0.350438 ;
  RECT 0.57881 0.04725 0.597185 0.216562 ;
  RECT 0.57881 0.216562 0.597185 0.332062 ;
  RECT 0.57881 0.332062 0.597185 0.350438 ;
  RECT 0.57881 0.350438 0.597185 0.441 ;
  RECT 0.662815 0.066872 0.681185 0.0853125 ;
  RECT 0.662815 0.0853125 0.681185 0.240187 ;
  RECT 0.662815 0.240187 0.681185 0.439688 ;
  RECT 0.681185 0.066872 0.876095 0.0853125 ;
  RECT 0.876095 0.066872 0.89447 0.0853125 ;
  RECT 0.876095 0.0853125 0.89447 0.240187 ;
  RECT 0.80325 0.258562 0.821625 0.418687 ;
  RECT 0.80325 0.418687 0.821625 0.437063 ;
  RECT 0.821625 0.418687 0.95681 0.437063 ;
  RECT 0.95681 0.04725 0.975185 0.086625 ;
  RECT 0.95681 0.086625 0.975185 0.258562 ;
  RECT 0.95681 0.258562 0.975185 0.418687 ;
  RECT 0.95681 0.418687 0.975185 0.437063 ;
  RECT 0.975185 0.086625 0.9765 0.258562 ;
  RECT 0.975185 0.258562 0.9765 0.418687 ;
  RECT 0.975185 0.418687 0.9765 0.437063 ;
  RECT 0.0315 0.055781 0.0525 0.0924655 ;
  RECT 0.0315 0.0924655 0.0525 0.110906 ;
  RECT 0.0315 0.372028 0.0525 0.397688 ;
  RECT 0.0315 0.397688 0.0525 0.450188 ;
  RECT 0.0525 0.0924655 0.0748125 0.110906 ;
  RECT 0.0525 0.372028 0.0748125 0.397688 ;
  RECT 0.0748125 0.0924655 0.093122 0.110906 ;
  RECT 0.0748125 0.110906 0.093122 0.372028 ;
  RECT 0.0748125 0.372028 0.093122 0.397688 ;
  RECT 0.242812 0.127312 0.261188 0.324188 ;
  RECT 0.326813 0.263813 0.345187 0.376688 ;
  RECT 0.345187 0.127312 0.366187 0.192937 ;
  RECT 0.483 0.169312 0.501375 0.287438 ;
  RECT 0.62081 0.179812 0.63919 0.379312 ;
  RECT 0.70481 0.114122 0.723185 0.208031 ;
  RECT 0.70481 0.301875 0.723185 0.408187 ;
  RECT 0.758625 0.108937 0.779625 0.450188 ;
  RECT 0.83081 0.114122 0.849185 0.208687 ;
      LAYER V1 ;
  RECT 0.0748125 0.347813 0.093122 0.366187 ;
  RECT 0.116812 0.137812 0.135187 0.156187 ;
  RECT 0.242812 0.137812 0.261188 0.156187 ;
  RECT 0.326813 0.347813 0.345187 0.366187 ;
  RECT 0.347813 0.137812 0.366187 0.156187 ;
  RECT 0.483 0.179812 0.501375 0.198187 ;
  RECT 0.62081 0.347813 0.63919 0.366187 ;
  RECT 0.70481 0.137812 0.723185 0.156187 ;
  RECT 0.70481 0.347813 0.723185 0.366187 ;
  RECT 0.83081 0.179812 0.849185 0.198187 ;
      LAYER M1 ;
  RECT 0.116812 0.04725 0.135187 0.456685 ;
  RECT 0.200812 0.04725 0.219187 0.456685 ;
  RECT 0.347813 0.408845 0.53412 0.446905 ;
  RECT 0.284813 0.066872 0.303187 0.0853125 ;
  RECT 0.284813 0.0853125 0.303187 0.287438 ;
  RECT 0.284813 0.287438 0.303187 0.439688 ;
  RECT 0.303187 0.066872 0.525 0.0853125 ;
  RECT 0.525 0.066872 0.543375 0.0853125 ;
  RECT 0.525 0.0853125 0.543375 0.287438 ;
  RECT 0.378 0.216562 0.396375 0.332062 ;
  RECT 0.378 0.332062 0.396375 0.350438 ;
  RECT 0.396375 0.332062 0.57881 0.350438 ;
  RECT 0.57881 0.04725 0.597185 0.216562 ;
  RECT 0.57881 0.216562 0.597185 0.332062 ;
  RECT 0.57881 0.332062 0.597185 0.350438 ;
  RECT 0.57881 0.350438 0.597185 0.441 ;
  RECT 0.662815 0.066872 0.681185 0.0853125 ;
  RECT 0.662815 0.0853125 0.681185 0.240187 ;
  RECT 0.662815 0.240187 0.681185 0.439688 ;
  RECT 0.681185 0.066872 0.876095 0.0853125 ;
  RECT 0.876095 0.066872 0.89447 0.0853125 ;
  RECT 0.876095 0.0853125 0.89447 0.240187 ;
  RECT 0.80325 0.258562 0.821625 0.418687 ;
  RECT 0.80325 0.418687 0.821625 0.437063 ;
  RECT 0.821625 0.418687 0.95681 0.437063 ;
  RECT 0.95681 0.04725 0.975185 0.086625 ;
  RECT 0.95681 0.086625 0.975185 0.258562 ;
  RECT 0.95681 0.258562 0.975185 0.418687 ;
  RECT 0.95681 0.418687 0.975185 0.437063 ;
  RECT 0.975185 0.086625 0.9765 0.258562 ;
  RECT 0.975185 0.258562 0.9765 0.418687 ;
  RECT 0.975185 0.418687 0.9765 0.437063 ;
  RECT 0.0315 0.055781 0.0525 0.0924655 ;
  RECT 0.0315 0.0924655 0.0525 0.110906 ;
  RECT 0.0315 0.372028 0.0525 0.397688 ;
  RECT 0.0315 0.397688 0.0525 0.450188 ;
  RECT 0.0525 0.0924655 0.0748125 0.110906 ;
  RECT 0.0525 0.372028 0.0748125 0.397688 ;
  RECT 0.0748125 0.0924655 0.093122 0.110906 ;
  RECT 0.0748125 0.110906 0.093122 0.372028 ;
  RECT 0.0748125 0.372028 0.093122 0.397688 ;
  RECT 0.242812 0.127312 0.261188 0.324188 ;
  RECT 0.326813 0.263813 0.345187 0.376688 ;
  RECT 0.345187 0.127312 0.366187 0.192937 ;
  RECT 0.483 0.169312 0.501375 0.287438 ;
  RECT 0.62081 0.179812 0.63919 0.379312 ;
  RECT 0.70481 0.114122 0.723185 0.208031 ;
  RECT 0.70481 0.301875 0.723185 0.408187 ;
  RECT 0.758625 0.108937 0.779625 0.450188 ;
  RECT 0.83081 0.114122 0.849185 0.208687 ;
  END
END DFFRNQ_X1

MACRO DFFSNQ_X1
  CLASS core ;
  FOREIGN DFFSNQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 1.092 BY 0.504 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.158812 0.177187 0.345187 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
  RECT 0.473813 0.179812 0.744125 0.198187 ;
  RECT 0.744125 0.179812 0.87019 0.198187 ;
    END
  END SN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.168 0.0511875 0.336 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 1.0395 0.042 1.0605 0.462 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.093122 0.522375 ;
  RECT 0.093122 0.485625 0.135187 0.522375 ;
  RECT 0.135187 0.485625 0.219187 0.522375 ;
  RECT 0.219187 0.485625 0.261188 0.522375 ;
  RECT 0.261188 0.485625 0.345187 0.522375 ;
  RECT 0.345187 0.485625 0.363563 0.522375 ;
  RECT 0.363563 0.485625 0.597185 0.522375 ;
  RECT 0.597185 0.485625 0.63919 0.522375 ;
  RECT 0.63919 0.485625 0.72581 0.522375 ;
  RECT 0.72581 0.485625 0.91212 0.522375 ;
  RECT 0.91212 0.485625 0.9765 0.522375 ;
  RECT 0.9765 0.485625 1.09856 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 1.09856 0.018375 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
  RECT 0.0958125 0.137812 0.744125 0.156187 ;
  RECT 0.0538125 0.347813 0.744125 0.366187 ;
      LAYER MINT1 ;
  RECT 0.0958125 0.137812 0.744125 0.156187 ;
  RECT 0.0538125 0.347813 0.744125 0.366187 ;
      LAYER M1 ;
  RECT 0.116812 0.04725 0.135187 0.456685 ;
  RECT 0.200812 0.04725 0.219187 0.456685 ;
  RECT 0.284813 0.0800625 0.303187 0.0984375 ;
  RECT 0.284813 0.0984375 0.303187 0.240187 ;
  RECT 0.284813 0.240187 0.303187 0.439688 ;
  RECT 0.303187 0.0800625 0.53675 0.0984375 ;
  RECT 0.53675 0.0800625 0.555185 0.0984375 ;
  RECT 0.53675 0.0984375 0.555185 0.240187 ;
  RECT 0.62081 0.179812 0.63919 0.376688 ;
  RECT 0.70481 0.127312 0.72581 0.213281 ;
  RECT 0.70481 0.257905 0.72581 0.389813 ;
  RECT 0.83081 0.122062 0.849185 0.208687 ;
  RECT 0.788815 0.258562 0.807185 0.376688 ;
  RECT 0.788815 0.376688 0.807185 0.395062 ;
  RECT 0.807185 0.376688 0.95681 0.395062 ;
  RECT 0.95681 0.04725 0.975185 0.086625 ;
  RECT 0.95681 0.086625 0.975185 0.258562 ;
  RECT 0.95681 0.258562 0.975185 0.376688 ;
  RECT 0.95681 0.376688 0.975185 0.395062 ;
  RECT 0.975185 0.086625 0.9765 0.258562 ;
  RECT 0.975185 0.258562 0.9765 0.376688 ;
  RECT 0.975185 0.376688 0.9765 0.395062 ;
  RECT 0.0295312 0.0538125 0.0315 0.0905625 ;
  RECT 0.0295312 0.0905625 0.0315 0.116156 ;
  RECT 0.0315 0.0538125 0.0525 0.0905625 ;
  RECT 0.0315 0.0905625 0.0525 0.116156 ;
  RECT 0.0315 0.372028 0.0525 0.397688 ;
  RECT 0.0315 0.397688 0.0525 0.450188 ;
  RECT 0.0525 0.0538125 0.054469 0.0905625 ;
  RECT 0.0525 0.0905625 0.054469 0.116156 ;
  RECT 0.0525 0.372028 0.054469 0.397688 ;
  RECT 0.054469 0.0905625 0.0748125 0.116156 ;
  RECT 0.054469 0.372028 0.0748125 0.397688 ;
  RECT 0.0748125 0.0905625 0.093122 0.116156 ;
  RECT 0.0748125 0.116156 0.093122 0.372028 ;
  RECT 0.0748125 0.372028 0.093122 0.397688 ;
  RECT 0.242812 0.127312 0.261188 0.324188 ;
  RECT 0.326813 0.263813 0.345187 0.387188 ;
  RECT 0.345187 0.127312 0.363563 0.200156 ;
  RECT 0.494812 0.169312 0.51319 0.240187 ;
  RECT 0.399 0.179812 0.417375 0.376688 ;
  RECT 0.399 0.376688 0.417375 0.395062 ;
  RECT 0.417375 0.376688 0.576185 0.395062 ;
  RECT 0.576185 0.376688 0.57881 0.395062 ;
  RECT 0.576185 0.395062 0.57881 0.450188 ;
  RECT 0.57881 0.063 0.597185 0.179812 ;
  RECT 0.57881 0.179812 0.597185 0.376688 ;
  RECT 0.57881 0.376688 0.597185 0.395062 ;
  RECT 0.57881 0.395062 0.597185 0.450188 ;
  RECT 0.662815 0.0748125 0.681185 0.093122 ;
  RECT 0.662815 0.093122 0.681185 0.240187 ;
  RECT 0.662815 0.240187 0.681185 0.441 ;
  RECT 0.681185 0.0748125 0.88725 0.093122 ;
  RECT 0.88725 0.0748125 0.90556 0.093122 ;
  RECT 0.88725 0.093122 0.90556 0.240187 ;
  RECT 0.72581 0.418687 0.91212 0.437063 ;
      LAYER V1 ;
  RECT 0.0748125 0.347813 0.093122 0.366187 ;
  RECT 0.116812 0.137812 0.135187 0.156187 ;
  RECT 0.242812 0.137812 0.261188 0.156187 ;
  RECT 0.326813 0.347813 0.345187 0.366187 ;
  RECT 0.345187 0.137812 0.363563 0.156187 ;
  RECT 0.494812 0.179812 0.51319 0.198187 ;
  RECT 0.62081 0.347813 0.63919 0.366187 ;
  RECT 0.70481 0.137812 0.723185 0.156187 ;
  RECT 0.70481 0.347813 0.723185 0.366187 ;
  RECT 0.83081 0.179812 0.849185 0.198187 ;
      LAYER M1 ;
  RECT 0.116812 0.04725 0.135187 0.456685 ;
  RECT 0.200812 0.04725 0.219187 0.456685 ;
  RECT 0.284813 0.0800625 0.303187 0.0984375 ;
  RECT 0.284813 0.0984375 0.303187 0.240187 ;
  RECT 0.284813 0.240187 0.303187 0.439688 ;
  RECT 0.303187 0.0800625 0.53675 0.0984375 ;
  RECT 0.53675 0.0800625 0.555185 0.0984375 ;
  RECT 0.53675 0.0984375 0.555185 0.240187 ;
  RECT 0.62081 0.179812 0.63919 0.376688 ;
  RECT 0.70481 0.127312 0.72581 0.213281 ;
  RECT 0.70481 0.257905 0.72581 0.389813 ;
  RECT 0.83081 0.122062 0.849185 0.208687 ;
  RECT 0.788815 0.258562 0.807185 0.376688 ;
  RECT 0.788815 0.376688 0.807185 0.395062 ;
  RECT 0.807185 0.376688 0.95681 0.395062 ;
  RECT 0.95681 0.04725 0.975185 0.086625 ;
  RECT 0.95681 0.086625 0.975185 0.258562 ;
  RECT 0.95681 0.258562 0.975185 0.376688 ;
  RECT 0.95681 0.376688 0.975185 0.395062 ;
  RECT 0.975185 0.086625 0.9765 0.258562 ;
  RECT 0.975185 0.258562 0.9765 0.376688 ;
  RECT 0.975185 0.376688 0.9765 0.395062 ;
  RECT 0.0295312 0.0538125 0.0315 0.0905625 ;
  RECT 0.0295312 0.0905625 0.0315 0.116156 ;
  RECT 0.0315 0.0538125 0.0525 0.0905625 ;
  RECT 0.0315 0.0905625 0.0525 0.116156 ;
  RECT 0.0315 0.372028 0.0525 0.397688 ;
  RECT 0.0315 0.397688 0.0525 0.450188 ;
  RECT 0.0525 0.0538125 0.054469 0.0905625 ;
  RECT 0.0525 0.0905625 0.054469 0.116156 ;
  RECT 0.0525 0.372028 0.054469 0.397688 ;
  RECT 0.054469 0.0905625 0.0748125 0.116156 ;
  RECT 0.054469 0.372028 0.0748125 0.397688 ;
  RECT 0.0748125 0.0905625 0.093122 0.116156 ;
  RECT 0.0748125 0.116156 0.093122 0.372028 ;
  RECT 0.0748125 0.372028 0.093122 0.397688 ;
  RECT 0.242812 0.127312 0.261188 0.324188 ;
  RECT 0.326813 0.263813 0.345187 0.387188 ;
  RECT 0.345187 0.127312 0.363563 0.200156 ;
  RECT 0.494812 0.169312 0.51319 0.240187 ;
  RECT 0.399 0.179812 0.417375 0.376688 ;
  RECT 0.399 0.376688 0.417375 0.395062 ;
  RECT 0.417375 0.376688 0.576185 0.395062 ;
  RECT 0.576185 0.376688 0.57881 0.395062 ;
  RECT 0.576185 0.395062 0.57881 0.450188 ;
  RECT 0.57881 0.063 0.597185 0.179812 ;
  RECT 0.57881 0.179812 0.597185 0.376688 ;
  RECT 0.57881 0.376688 0.597185 0.395062 ;
  RECT 0.57881 0.395062 0.597185 0.450188 ;
  RECT 0.662815 0.0748125 0.681185 0.093122 ;
  RECT 0.662815 0.093122 0.681185 0.240187 ;
  RECT 0.662815 0.240187 0.681185 0.441 ;
  RECT 0.681185 0.0748125 0.88725 0.093122 ;
  RECT 0.88725 0.0748125 0.90556 0.093122 ;
  RECT 0.88725 0.093122 0.90556 0.240187 ;
  RECT 0.72581 0.418687 0.91212 0.437063 ;
  END
END DFFSNQ_X1

MACRO INV_X1
  CLASS core ;
  FOREIGN INV_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.126 BY 0.504 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.126 0.0511875 0.378 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.0748125 0.093122 0.42 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.132562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.132562 0.018375 ;
    END
  END VSS
END INV_X1

MACRO INV_X2
  CLASS core ;
  FOREIGN INV_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.126 BY 0.504 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.025 0.126 0.038 0.378   ; 
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.056 0.085 0.070 0.378   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.005 0.486 0.131 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.005 -0.018 0.131 0.018   ; 
    END
  END VSS
END INV_X2

MACRO INV_X4
  CLASS core ;
  FOREIGN INV_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.126 BY 0.504 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.016 0.168 0.026 0.241   ; 
  RECT 0.016 0.241 0.026 0.260   ; 
  RECT 0.016 0.260 0.026 0.336   ; 
  RECT 0.026 0.241 0.078 0.260   ; 
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.013 0.093 0.019 0.131   ; 
  RECT 0.019 0.093 0.100 0.131   ; 
  RECT 0.019 0.373 0.100 0.411   ; 
  RECT 0.100 0.093 0.110 0.131   ; 
  RECT 0.100 0.131 0.110 0.373   ; 
  RECT 0.100 0.373 0.110 0.411   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.003 0.486 0.129 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.003 -0.018 0.129 0.018   ; 
    END
  END VSS
END INV_X4

MACRO INV_X8
  CLASS core ;
  FOREIGN INV_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.126 BY 0.504 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.022 0.127 0.028 0.260   ; 
  RECT 0.022 0.260 0.028 0.299   ; 
  RECT 0.022 0.299 0.028 0.378   ; 
  RECT 0.028 0.260 0.091 0.299   ; 
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.008 0.414 0.011 0.432   ; 
  RECT 0.011 0.072 0.110 0.091   ; 
  RECT 0.011 0.414 0.110 0.432   ; 
  RECT 0.110 0.072 0.117 0.091   ; 
  RECT 0.110 0.091 0.117 0.414   ; 
  RECT 0.110 0.414 0.117 0.432   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.002 0.486 0.128 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.002 -0.018 0.128 0.018   ; 
    END
  END VSS
END INV_X8

MACRO INV_X12
  CLASS core ;
  FOREIGN INV_X12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.168 BY 0.504 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.021 0.126 0.027 0.241   ; 
  RECT 0.021 0.241 0.027 0.260   ; 
  RECT 0.021 0.260 0.027 0.378   ; 
  RECT 0.027 0.241 0.129 0.260   ; 
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.010 0.067 0.152 0.085   ; 
  RECT 0.010 0.417 0.152 0.438   ; 
  RECT 0.152 0.067 0.160 0.085   ; 
  RECT 0.152 0.085 0.160 0.417   ; 
  RECT 0.152 0.417 0.160 0.438   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.002 0.486 0.170 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.002 -0.018 0.170 0.018   ; 
    END
  END VSS
END INV_X12

MACRO INV_X16
  CLASS core ;
  FOREIGN INV_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.168 BY 0.504 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.007 0.168 0.011 0.243   ; 
  RECT 0.007 0.243 0.011 0.261   ; 
  RECT 0.007 0.261 0.011 0.369   ; 
  RECT 0.011 0.243 0.137 0.261   ; 
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.001 0.486 0.156 0.522   ; 
  RECT 0.156 0.486 0.169 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.001 -0.018 0.169 0.018   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.008 0.066 0.151 0.087   ; 
  RECT 0.008 0.408 0.151 0.447   ; 
  RECT 0.151 0.066 0.156 0.087   ; 
  RECT 0.151 0.087 0.156 0.408   ; 
  RECT 0.151 0.408 0.156 0.447   ; 
      LAYER M1 ;
  RECT 0.008 0.066 0.151 0.087   ; 
  RECT 0.008 0.408 0.151 0.447   ; 
  RECT 0.151 0.066 0.156 0.087   ; 
  RECT 0.151 0.087 0.156 0.408   ; 
  RECT 0.151 0.408 0.156 0.447   ; 
  END
END INV_X16

MACRO LHQ_X1
  CLASS core ;
  FOREIGN LHQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.588 BY 0.504 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.105 0.177187 0.336 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.168 0.0511875 0.336 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.53675 0.0853125 0.555185 0.418687 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.51319 0.522375 ;
  RECT 0.51319 0.485625 0.59456 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.59456 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0315 0.364875 0.0328125 0.38325 ;
  RECT 0.0315 0.38325 0.0328125 0.462 ;
  RECT 0.0328125 0.042 0.0511875 0.060375 ;
  RECT 0.0328125 0.060375 0.0511875 0.12075 ;
  RECT 0.0328125 0.12075 0.0511875 0.139125 ;
  RECT 0.0328125 0.364875 0.0511875 0.38325 ;
  RECT 0.0328125 0.38325 0.0511875 0.462 ;
  RECT 0.0511875 0.042 0.0525 0.060375 ;
  RECT 0.0511875 0.12075 0.0525 0.139125 ;
  RECT 0.0511875 0.364875 0.0525 0.38325 ;
  RECT 0.0511875 0.38325 0.0525 0.462 ;
  RECT 0.0525 0.042 0.0748125 0.060375 ;
  RECT 0.0525 0.12075 0.0748125 0.139125 ;
  RECT 0.0525 0.364875 0.0748125 0.38325 ;
  RECT 0.0748125 0.042 0.093122 0.060375 ;
  RECT 0.0748125 0.12075 0.093122 0.139125 ;
  RECT 0.0748125 0.139125 0.093122 0.211312 ;
  RECT 0.0748125 0.211312 0.093122 0.229687 ;
  RECT 0.0748125 0.229687 0.093122 0.271688 ;
  RECT 0.0748125 0.271688 0.093122 0.364875 ;
  RECT 0.0748125 0.364875 0.093122 0.38325 ;
  RECT 0.093122 0.042 0.212625 0.060375 ;
  RECT 0.212625 0.042 0.231 0.060375 ;
  RECT 0.212625 0.060375 0.231 0.12075 ;
  RECT 0.212625 0.12075 0.231 0.139125 ;
  RECT 0.212625 0.139125 0.231 0.211312 ;
  RECT 0.212625 0.211312 0.231 0.229687 ;
  RECT 0.231 0.211312 0.242812 0.229687 ;
  RECT 0.242812 0.211312 0.261188 0.229687 ;
  RECT 0.242812 0.229687 0.261188 0.271688 ;
  RECT 0.347813 0.0748125 0.366187 0.093122 ;
  RECT 0.347813 0.093122 0.366187 0.324188 ;
  RECT 0.366187 0.0748125 0.452748 0.093122 ;
  RECT 0.452748 0.0748125 0.471187 0.093122 ;
  RECT 0.452748 0.093122 0.471187 0.324188 ;
  RECT 0.452748 0.324188 0.471187 0.389155 ;
  RECT 0.116812 0.08925 0.135187 0.301875 ;
  RECT 0.116812 0.301875 0.135187 0.364875 ;
  RECT 0.116812 0.364875 0.135187 0.38325 ;
  RECT 0.135187 0.364875 0.200812 0.38325 ;
  RECT 0.200812 0.301875 0.223125 0.364875 ;
  RECT 0.200812 0.364875 0.223125 0.38325 ;
  RECT 0.179812 0.418687 0.254625 0.437063 ;
  RECT 0.254625 0.0748125 0.305812 0.113466 ;
  RECT 0.254625 0.418687 0.305812 0.437063 ;
  RECT 0.305812 0.0748125 0.324188 0.113466 ;
  RECT 0.305812 0.113466 0.324188 0.200812 ;
  RECT 0.305812 0.200812 0.324188 0.41803 ;
  RECT 0.305812 0.41803 0.324188 0.418687 ;
  RECT 0.305812 0.418687 0.324188 0.437063 ;
  RECT 0.324188 0.41803 0.494812 0.418687 ;
  RECT 0.324188 0.418687 0.494812 0.437063 ;
  RECT 0.494812 0.200812 0.51319 0.41803 ;
  RECT 0.494812 0.41803 0.51319 0.418687 ;
  RECT 0.494812 0.418687 0.51319 0.437063 ;
      LAYER M1 ;
  RECT 0.0315 0.364875 0.0328125 0.38325 ;
  RECT 0.0315 0.38325 0.0328125 0.462 ;
  RECT 0.0328125 0.042 0.0511875 0.060375 ;
  RECT 0.0328125 0.060375 0.0511875 0.12075 ;
  RECT 0.0328125 0.12075 0.0511875 0.139125 ;
  RECT 0.0328125 0.364875 0.0511875 0.38325 ;
  RECT 0.0328125 0.38325 0.0511875 0.462 ;
  RECT 0.0511875 0.042 0.0525 0.060375 ;
  RECT 0.0511875 0.12075 0.0525 0.139125 ;
  RECT 0.0511875 0.364875 0.0525 0.38325 ;
  RECT 0.0511875 0.38325 0.0525 0.462 ;
  RECT 0.0525 0.042 0.0748125 0.060375 ;
  RECT 0.0525 0.12075 0.0748125 0.139125 ;
  RECT 0.0525 0.364875 0.0748125 0.38325 ;
  RECT 0.0748125 0.042 0.093122 0.060375 ;
  RECT 0.0748125 0.12075 0.093122 0.139125 ;
  RECT 0.0748125 0.139125 0.093122 0.211312 ;
  RECT 0.0748125 0.211312 0.093122 0.229687 ;
  RECT 0.0748125 0.229687 0.093122 0.271688 ;
  RECT 0.0748125 0.271688 0.093122 0.364875 ;
  RECT 0.0748125 0.364875 0.093122 0.38325 ;
  RECT 0.093122 0.042 0.212625 0.060375 ;
  RECT 0.212625 0.042 0.231 0.060375 ;
  RECT 0.212625 0.060375 0.231 0.12075 ;
  RECT 0.212625 0.12075 0.231 0.139125 ;
  RECT 0.212625 0.139125 0.231 0.211312 ;
  RECT 0.212625 0.211312 0.231 0.229687 ;
  RECT 0.231 0.211312 0.242812 0.229687 ;
  RECT 0.242812 0.211312 0.261188 0.229687 ;
  RECT 0.242812 0.229687 0.261188 0.271688 ;
  RECT 0.347813 0.0748125 0.366187 0.093122 ;
  RECT 0.347813 0.093122 0.366187 0.324188 ;
  RECT 0.366187 0.0748125 0.452748 0.093122 ;
  RECT 0.452748 0.0748125 0.471187 0.093122 ;
  RECT 0.452748 0.093122 0.471187 0.324188 ;
  RECT 0.452748 0.324188 0.471187 0.389155 ;
  RECT 0.116812 0.08925 0.135187 0.301875 ;
  RECT 0.116812 0.301875 0.135187 0.364875 ;
  RECT 0.116812 0.364875 0.135187 0.38325 ;
  RECT 0.135187 0.364875 0.200812 0.38325 ;
  RECT 0.200812 0.301875 0.223125 0.364875 ;
  RECT 0.200812 0.364875 0.223125 0.38325 ;
  RECT 0.179812 0.418687 0.254625 0.437063 ;
  RECT 0.254625 0.0748125 0.305812 0.113466 ;
  RECT 0.254625 0.418687 0.305812 0.437063 ;
  RECT 0.305812 0.0748125 0.324188 0.113466 ;
  RECT 0.305812 0.113466 0.324188 0.200812 ;
  RECT 0.305812 0.200812 0.324188 0.41803 ;
  RECT 0.305812 0.41803 0.324188 0.418687 ;
  RECT 0.305812 0.418687 0.324188 0.437063 ;
  RECT 0.324188 0.41803 0.494812 0.418687 ;
  RECT 0.324188 0.418687 0.494812 0.437063 ;
  RECT 0.494812 0.200812 0.51319 0.41803 ;
  RECT 0.494812 0.41803 0.51319 0.418687 ;
  RECT 0.494812 0.418687 0.51319 0.437063 ;
  END
END LHQ_X1

MACRO MUX2_X1
  CLASS core ;
  FOREIGN MUX2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.546 BY 0.504 ;
  PIN I0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.368812 0.158812 0.387188 0.345187 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.168 0.093122 0.294 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
  RECT 0.0774375 0.431812 0.258562 0.450188 ;
      LAYER V1 ;
  RECT 0.0984375 0.431812 0.135187 0.450188 ;
      LAYER M1 ;
  RECT 0.0177187 0.158812 0.0360938 0.431812 ;
  RECT 0.0177187 0.431812 0.0360938 0.450188 ;
  RECT 0.0360938 0.431812 0.145687 0.450188 ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.452748 0.126 0.471187 0.418687 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.303187 0.522375 ;
  RECT 0.303187 0.485625 0.345187 0.522375 ;
  RECT 0.345187 0.485625 0.51319 0.522375 ;
  RECT 0.51319 0.485625 0.55256 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.55256 0.018375 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
  RECT 0.179812 0.221812 0.366187 0.240187 ;
      LAYER MINT1 ;
  RECT 0.179812 0.221812 0.366187 0.240187 ;
      LAYER M1 ;
  RECT 0.0525 0.106312 0.064969 0.124687 ;
  RECT 0.064969 0.106312 0.103031 0.124687 ;
  RECT 0.064969 0.322875 0.103031 0.34125 ;
  RECT 0.064969 0.34125 0.103031 0.378 ;
  RECT 0.103031 0.106312 0.200812 0.124687 ;
  RECT 0.103031 0.322875 0.200812 0.34125 ;
  RECT 0.200812 0.106312 0.219187 0.124687 ;
  RECT 0.200812 0.124687 0.219187 0.322875 ;
  RECT 0.200812 0.322875 0.219187 0.34125 ;
  RECT 0.190312 0.431812 0.284813 0.462 ;
  RECT 0.284813 0.200812 0.303187 0.431812 ;
  RECT 0.284813 0.431812 0.303187 0.462 ;
  RECT 0.326813 0.179812 0.345187 0.280875 ;
  RECT 0.242812 0.057028 0.261188 0.0958125 ;
  RECT 0.242812 0.0958125 0.261188 0.324188 ;
  RECT 0.242812 0.324188 0.261188 0.402938 ;
  RECT 0.261188 0.057028 0.494812 0.0958125 ;
  RECT 0.494812 0.057028 0.51319 0.0958125 ;
  RECT 0.494812 0.0958125 0.51319 0.324188 ;
      LAYER V1 ;
  RECT 0.200812 0.221812 0.219187 0.240187 ;
  RECT 0.200812 0.431812 0.237562 0.450188 ;
  RECT 0.326813 0.221812 0.345187 0.240187 ;
      LAYER M1 ;
  RECT 0.0525 0.106312 0.064969 0.124687 ;
  RECT 0.064969 0.106312 0.103031 0.124687 ;
  RECT 0.064969 0.322875 0.103031 0.34125 ;
  RECT 0.064969 0.34125 0.103031 0.378 ;
  RECT 0.103031 0.106312 0.200812 0.124687 ;
  RECT 0.103031 0.322875 0.200812 0.34125 ;
  RECT 0.200812 0.106312 0.219187 0.124687 ;
  RECT 0.200812 0.124687 0.219187 0.322875 ;
  RECT 0.200812 0.322875 0.219187 0.34125 ;
  RECT 0.190312 0.431812 0.284813 0.462 ;
  RECT 0.284813 0.200812 0.303187 0.431812 ;
  RECT 0.284813 0.431812 0.303187 0.462 ;
  RECT 0.326813 0.179812 0.345187 0.280875 ;
  RECT 0.242812 0.057028 0.261188 0.0958125 ;
  RECT 0.242812 0.0958125 0.261188 0.324188 ;
  RECT 0.242812 0.324188 0.261188 0.402938 ;
  RECT 0.261188 0.057028 0.494812 0.0958125 ;
  RECT 0.494812 0.057028 0.51319 0.0958125 ;
  RECT 0.494812 0.0958125 0.51319 0.324188 ;
  END
END MUX2_X1

MACRO NAND2_X1
  CLASS core ;
  FOREIGN NAND2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.168 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.168 0.135187 0.376688 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.168 0.0511875 0.376688 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.0872815 0.093122 0.126 ;
  RECT 0.0748125 0.126 0.093122 0.418687 ;
  RECT 0.093122 0.0872815 0.1155 0.126 ;
  RECT 0.1155 0.042 0.1365 0.0872815 ;
  RECT 0.1155 0.0872815 0.1365 0.126 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.174562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.174562 0.018375 ;
    END
  END VSS
END NAND2_X1

MACRO NAND2_X2
  CLASS core ;
  FOREIGN NAND2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.168 BY 0.504 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.078 0.148 0.090 0.363   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.022 0.180 0.034 0.444   ; 
  RECT 0.022 0.444 0.034 0.462   ; 
  RECT 0.034 0.444 0.134 0.462   ; 
  RECT 0.134 0.180 0.146 0.444   ; 
  RECT 0.134 0.444 0.146 0.462   ; 
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.050 0.081 0.062 0.119   ; 
  RECT 0.050 0.119 0.062 0.278   ; 
  RECT 0.050 0.278 0.062 0.392   ; 
  RECT 0.050 0.392 0.062 0.420   ; 
  RECT 0.062 0.081 0.106 0.119   ; 
  RECT 0.062 0.392 0.106 0.420   ; 
  RECT 0.106 0.081 0.118 0.119   ; 
  RECT 0.106 0.278 0.118 0.392   ; 
  RECT 0.106 0.392 0.118 0.420   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.004 0.486 0.172 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.004 -0.018 0.172 0.018   ; 
    END
  END VSS
END NAND2_X2

MACRO NAND3_X1
  CLASS core ;
  FOREIGN NAND3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.252 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.21 0.177187 0.294 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.167344 0.135187 0.336 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.141094 0.0511875 0.376688 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.0538125 0.093122 0.0721875 ;
  RECT 0.0748125 0.0721875 0.093122 0.168 ;
  RECT 0.0748125 0.168 0.093122 0.336 ;
  RECT 0.0748125 0.336 0.093122 0.443625 ;
  RECT 0.0748125 0.443625 0.093122 0.462 ;
  RECT 0.093122 0.0538125 0.158812 0.0721875 ;
  RECT 0.093122 0.443625 0.158812 0.462 ;
  RECT 0.158812 0.042 0.1995 0.0538125 ;
  RECT 0.158812 0.0538125 0.1995 0.0721875 ;
  RECT 0.158812 0.443625 0.1995 0.462 ;
  RECT 0.1995 0.042 0.200812 0.0538125 ;
  RECT 0.1995 0.0538125 0.200812 0.0721875 ;
  RECT 0.1995 0.0721875 0.200812 0.168 ;
  RECT 0.1995 0.443625 0.200812 0.462 ;
  RECT 0.200812 0.042 0.219187 0.0538125 ;
  RECT 0.200812 0.0538125 0.219187 0.0721875 ;
  RECT 0.200812 0.0721875 0.219187 0.168 ;
  RECT 0.200812 0.336 0.219187 0.443625 ;
  RECT 0.200812 0.443625 0.219187 0.462 ;
  RECT 0.219187 0.042 0.2205 0.0538125 ;
  RECT 0.219187 0.0538125 0.2205 0.0721875 ;
  RECT 0.219187 0.0721875 0.2205 0.168 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.258562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.258562 0.018375 ;
    END
  END VSS
END NAND3_X1

MACRO NAND3_X2
  CLASS core ;
  FOREIGN NAND3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.252 BY 0.504 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.218 0.210 0.230 0.336   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.132 0.163 0.148 0.336   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.050 0.168 0.062 0.336   ; 
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.012 0.373 0.160 0.411   ; 
  RECT 0.160 0.373 0.190 0.411   ; 
  RECT 0.190 0.122 0.202 0.373   ; 
  RECT 0.190 0.373 0.202 0.411   ; 
  RECT 0.202 0.373 0.216 0.411   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.004 0.486 0.160 0.522   ; 
  RECT 0.160 0.486 0.230 0.522   ; 
  RECT 0.230 0.486 0.256 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.004 -0.018 0.256 0.018   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.092 0.073 0.218 0.092   ; 
  RECT 0.218 0.073 0.230 0.092   ; 
  RECT 0.218 0.092 0.230 0.148   ; 
  RECT 0.022 0.116 0.160 0.137   ; 
      LAYER M1 ;
  RECT 0.092 0.073 0.218 0.092   ; 
  RECT 0.218 0.073 0.230 0.092   ; 
  RECT 0.218 0.092 0.230 0.148   ; 
  RECT 0.022 0.116 0.160 0.137   ; 
  END
END NAND3_X2

MACRO NAND4_X1
  CLASS core ;
  FOREIGN NAND4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.294 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.242812 0.168 0.261188 0.376688 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.158812 0.177187 0.336 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.127312 0.135187 0.294 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.127312 0.0511875 0.376688 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.336 0.093122 0.42328 ;
  RECT 0.0748125 0.42328 0.093122 0.462 ;
  RECT 0.093122 0.42328 0.200812 0.462 ;
  RECT 0.200812 0.107625 0.219187 0.126 ;
  RECT 0.200812 0.126 0.219187 0.336 ;
  RECT 0.200812 0.336 0.219187 0.42328 ;
  RECT 0.200812 0.42328 0.219187 0.462 ;
  RECT 0.219187 0.107625 0.239531 0.126 ;
  RECT 0.239531 0.042 0.26447 0.107625 ;
  RECT 0.239531 0.107625 0.26447 0.126 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.300563 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.300563 0.018375 ;
    END
  END VSS
END NAND4_X1

MACRO NAND4_X2
  CLASS core ;
  FOREIGN NAND4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.294 BY 0.504 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.233 0.235 0.248 0.336   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.155 0.223 0.166 0.345   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.074 0.159 0.086 0.336   ; 
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.021 0.169 0.033 0.336   ; 
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.047 0.364 0.060 0.378   ; 
  RECT 0.047 0.378 0.060 0.419   ; 
  RECT 0.047 0.419 0.060 0.437   ; 
  RECT 0.060 0.419 0.181 0.437   ; 
  RECT 0.181 0.193 0.193 0.211   ; 
  RECT 0.181 0.211 0.193 0.360   ; 
  RECT 0.181 0.360 0.193 0.364   ; 
  RECT 0.181 0.364 0.193 0.378   ; 
  RECT 0.181 0.419 0.193 0.437   ; 
  RECT 0.193 0.193 0.235 0.211   ; 
  RECT 0.193 0.360 0.235 0.364   ; 
  RECT 0.193 0.364 0.235 0.378   ; 
  RECT 0.193 0.419 0.235 0.437   ; 
  RECT 0.235 0.193 0.246 0.211   ; 
  RECT 0.235 0.360 0.246 0.364   ; 
  RECT 0.235 0.364 0.246 0.378   ; 
  RECT 0.235 0.378 0.246 0.419   ; 
  RECT 0.235 0.419 0.246 0.437   ; 
  RECT 0.246 0.193 0.273 0.211   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.004 0.486 0.274 0.522   ; 
  RECT 0.274 0.486 0.298 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.004 -0.018 0.298 0.018   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.020 0.067 0.033 0.085   ; 
  RECT 0.020 0.085 0.033 0.140   ; 
  RECT 0.033 0.067 0.180 0.085   ; 
  RECT 0.114 0.151 0.261 0.169   ; 
  RECT 0.261 0.042 0.274 0.151   ; 
  RECT 0.261 0.151 0.274 0.169   ; 
  RECT 0.061 0.109 0.206 0.127   ; 
      LAYER M1 ;
  RECT 0.020 0.067 0.033 0.085   ; 
  RECT 0.020 0.085 0.033 0.140   ; 
  RECT 0.033 0.067 0.180 0.085   ; 
  RECT 0.114 0.151 0.261 0.169   ; 
  RECT 0.261 0.042 0.274 0.151   ; 
  RECT 0.261 0.151 0.274 0.169   ; 
  RECT 0.061 0.109 0.206 0.127   ; 
  END
END NAND4_X2

MACRO NOR2_X1
  CLASS core ;
  FOREIGN NOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.168 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.127312 0.135187 0.336 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.127312 0.0511875 0.336 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.0853125 0.093122 0.378 ;
  RECT 0.0748125 0.378 0.093122 0.41672 ;
  RECT 0.093122 0.378 0.1155 0.41672 ;
  RECT 0.1155 0.378 0.1365 0.41672 ;
  RECT 0.1155 0.41672 0.1365 0.462 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.174562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.174562 0.018375 ;
    END
  END VSS
END NOR2_X1

MACRO NOR2_X2
  CLASS core ;
  FOREIGN NOR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.168 BY 0.504 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.078 0.141 0.090 0.336   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.022 0.042 0.034 0.060   ; 
  RECT 0.022 0.060 0.034 0.324   ; 
  RECT 0.034 0.042 0.134 0.060   ; 
  RECT 0.134 0.042 0.146 0.060   ; 
  RECT 0.134 0.060 0.146 0.324   ; 
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.050 0.084 0.062 0.102   ; 
  RECT 0.050 0.102 0.062 0.226   ; 
  RECT 0.050 0.226 0.062 0.365   ; 
  RECT 0.050 0.365 0.062 0.383   ; 
  RECT 0.062 0.084 0.077 0.102   ; 
  RECT 0.062 0.365 0.077 0.383   ; 
  RECT 0.077 0.084 0.091 0.102   ; 
  RECT 0.077 0.365 0.091 0.383   ; 
  RECT 0.077 0.383 0.091 0.420   ; 
  RECT 0.091 0.084 0.106 0.102   ; 
  RECT 0.106 0.084 0.118 0.102   ; 
  RECT 0.106 0.102 0.118 0.226   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.004 0.486 0.172 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.004 -0.018 0.172 0.018   ; 
    END
  END VSS
END NOR2_X2

MACRO NOR3_X1
  CLASS core ;
  FOREIGN NOR3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.252 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.21 0.177187 0.294 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.127312 0.135187 0.362905 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.127312 0.0511875 0.362905 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.042 0.093122 0.060375 ;
  RECT 0.0748125 0.060375 0.093122 0.168 ;
  RECT 0.0748125 0.168 0.093122 0.336 ;
  RECT 0.0748125 0.336 0.093122 0.402938 ;
  RECT 0.0748125 0.402938 0.093122 0.421312 ;
  RECT 0.093122 0.042 0.198844 0.060375 ;
  RECT 0.093122 0.402938 0.198844 0.421312 ;
  RECT 0.198844 0.042 0.1995 0.060375 ;
  RECT 0.198844 0.060375 0.1995 0.168 ;
  RECT 0.198844 0.402938 0.1995 0.421312 ;
  RECT 0.1995 0.042 0.2205 0.060375 ;
  RECT 0.1995 0.060375 0.2205 0.168 ;
  RECT 0.1995 0.336 0.2205 0.402938 ;
  RECT 0.1995 0.402938 0.2205 0.421312 ;
  RECT 0.1995 0.421312 0.2205 0.462 ;
  RECT 0.2205 0.042 0.221156 0.060375 ;
  RECT 0.2205 0.060375 0.221156 0.168 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.258562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.258562 0.018375 ;
    END
  END VSS
END NOR3_X1

MACRO NOR3_X2
  CLASS core ;
  FOREIGN NOR3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.252 BY 0.504 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.218 0.168 0.230 0.294   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.134 0.168 0.146 0.337   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.022 0.168 0.034 0.341   ; 
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.038 0.101 0.190 0.139   ; 
  RECT 0.190 0.101 0.202 0.139   ; 
  RECT 0.190 0.139 0.202 0.378   ; 
  RECT 0.202 0.101 0.214 0.139   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.004 0.486 0.230 0.522   ; 
  RECT 0.230 0.486 0.256 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.004 -0.018 0.256 0.018   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.092 0.411 0.218 0.430   ; 
  RECT 0.218 0.339 0.230 0.411   ; 
  RECT 0.218 0.411 0.230 0.430   ; 
  RECT 0.038 0.366 0.166 0.388   ; 
      LAYER M1 ;
  RECT 0.092 0.411 0.218 0.430   ; 
  RECT 0.218 0.339 0.230 0.411   ; 
  RECT 0.218 0.411 0.230 0.430   ; 
  RECT 0.038 0.366 0.166 0.388   ; 
  END
END NOR3_X2

MACRO NOR4_X1
  CLASS core ;
  FOREIGN NOR4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.294 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.242812 0.127312 0.261188 0.336 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.127312 0.177187 0.336 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.168 0.135187 0.376688 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.127312 0.0511875 0.376688 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.042 0.093122 0.066872 ;
  RECT 0.0748125 0.066872 0.093122 0.141094 ;
  RECT 0.093122 0.042 0.200812 0.066872 ;
  RECT 0.200812 0.042 0.219187 0.066872 ;
  RECT 0.200812 0.066872 0.219187 0.141094 ;
  RECT 0.200812 0.141094 0.219187 0.378 ;
  RECT 0.200812 0.378 0.219187 0.396375 ;
  RECT 0.219187 0.378 0.239531 0.396375 ;
  RECT 0.239531 0.378 0.26447 0.396375 ;
  RECT 0.239531 0.396375 0.26447 0.462 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.300563 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.300563 0.018375 ;
    END
  END VSS
END NOR4_X1

MACRO NOR4_X2
  CLASS core ;
  FOREIGN NOR4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.294 BY 0.504 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.233 0.168 0.248 0.266   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.155 0.159 0.166 0.287   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.101 0.159 0.113 0.345   ; 
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.074 0.168 0.086 0.339   ; 
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.047 0.067 0.060 0.085   ; 
  RECT 0.047 0.085 0.060 0.126   ; 
  RECT 0.047 0.126 0.060 0.140   ; 
  RECT 0.060 0.067 0.181 0.085   ; 
  RECT 0.181 0.067 0.193 0.085   ; 
  RECT 0.181 0.126 0.193 0.140   ; 
  RECT 0.181 0.140 0.193 0.144   ; 
  RECT 0.181 0.144 0.193 0.290   ; 
  RECT 0.181 0.290 0.193 0.308   ; 
  RECT 0.193 0.067 0.235 0.085   ; 
  RECT 0.193 0.126 0.235 0.140   ; 
  RECT 0.193 0.140 0.235 0.144   ; 
  RECT 0.193 0.290 0.235 0.308   ; 
  RECT 0.235 0.067 0.246 0.085   ; 
  RECT 0.235 0.085 0.246 0.126   ; 
  RECT 0.235 0.126 0.246 0.140   ; 
  RECT 0.235 0.140 0.246 0.144   ; 
  RECT 0.235 0.290 0.246 0.308   ; 
  RECT 0.246 0.290 0.277 0.308   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.004 0.486 0.180 0.522   ; 
  RECT 0.180 0.486 0.206 0.522   ; 
  RECT 0.206 0.486 0.274 0.522   ; 
  RECT 0.274 0.486 0.298 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.004 -0.018 0.298 0.018   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.088 0.374 0.206 0.395   ; 
  RECT 0.020 0.364 0.033 0.419   ; 
  RECT 0.020 0.419 0.033 0.437   ; 
  RECT 0.033 0.419 0.180 0.437   ; 
  RECT 0.141 0.332 0.261 0.350   ; 
  RECT 0.261 0.332 0.274 0.350   ; 
  RECT 0.261 0.350 0.274 0.450   ; 
      LAYER M1 ;
  RECT 0.088 0.374 0.206 0.395   ; 
  RECT 0.020 0.364 0.033 0.419   ; 
  RECT 0.020 0.419 0.033 0.437   ; 
  RECT 0.033 0.419 0.180 0.437   ; 
  RECT 0.141 0.332 0.261 0.350   ; 
  RECT 0.261 0.332 0.274 0.350   ; 
  RECT 0.261 0.350 0.274 0.450   ; 
  END
END NOR4_X2


MACRO OAI21_X1
  CLASS core ;
  FOREIGN OAI21_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.252 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.168 0.135187 0.378 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.168 0.0511875 0.416063 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.200812 0.168 0.219187 0.378 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.168 0.093122 0.417375 ;
  RECT 0.0748125 0.417375 0.093122 0.438375 ;
  RECT 0.093122 0.417375 0.195562 0.438375 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.195562 0.522375 ;
  RECT 0.195562 0.485625 0.258562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.258562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0328125 0.0479062 0.0511875 0.101719 ;
  RECT 0.0328125 0.101719 0.0511875 0.122719 ;
  RECT 0.0511875 0.101719 0.195562 0.122719 ;
      LAYER M1 ;
  RECT 0.0328125 0.0479062 0.0511875 0.101719 ;
  RECT 0.0328125 0.101719 0.0511875 0.122719 ;
  RECT 0.0511875 0.101719 0.195562 0.122719 ;
  END
END OAI21_X1

MACRO OAI21_X2
  CLASS core ;
  FOREIGN OAI21_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.252 BY 0.504 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.160 0.210 0.176 0.294   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.106 0.159 0.118 0.186   ; 
  RECT 0.106 0.186 0.118 0.329   ; 
  RECT 0.106 0.329 0.118 0.348   ; 
  RECT 0.118 0.329 0.218 0.348   ; 
  RECT 0.218 0.186 0.230 0.329   ; 
  RECT 0.218 0.329 0.230 0.348   ; 
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.050 0.168 0.062 0.345   ; 
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.013 0.374 0.078 0.395   ; 
  RECT 0.078 0.109 0.090 0.127   ; 
  RECT 0.078 0.127 0.090 0.182   ; 
  RECT 0.078 0.182 0.090 0.374   ; 
  RECT 0.078 0.374 0.090 0.395   ; 
  RECT 0.090 0.109 0.186 0.127   ; 
  RECT 0.090 0.374 0.186 0.395   ; 
  RECT 0.186 0.109 0.190 0.127   ; 
  RECT 0.190 0.109 0.202 0.127   ; 
  RECT 0.190 0.127 0.202 0.182   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.004 0.486 0.234 0.522   ; 
  RECT 0.234 0.486 0.256 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.004 -0.018 0.256 0.018   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.021 0.067 0.035 0.085   ; 
  RECT 0.021 0.085 0.035 0.140   ; 
  RECT 0.035 0.067 0.218 0.085   ; 
  RECT 0.218 0.067 0.230 0.085   ; 
  RECT 0.218 0.085 0.230 0.140   ; 
  RECT 0.218 0.140 0.230 0.141   ; 
  RECT 0.064 0.419 0.234 0.437   ; 
      LAYER M1 ;
  RECT 0.021 0.067 0.035 0.085   ; 
  RECT 0.021 0.085 0.035 0.140   ; 
  RECT 0.035 0.067 0.218 0.085   ; 
  RECT 0.218 0.067 0.230 0.085   ; 
  RECT 0.218 0.085 0.230 0.140   ; 
  RECT 0.218 0.140 0.230 0.141   ; 
  RECT 0.064 0.419 0.234 0.437   ; 
  END
END OAI21_X2

MACRO OAI22_X1
  CLASS core ;
  FOREIGN OAI22_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.294 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.130594 0.177187 0.378 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.242812 0.183094 0.261188 0.378 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.126 0.135187 0.336 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0315 0.126 0.0525 0.378 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0924655 0.418687 0.200812 0.437063 ;
  RECT 0.200812 0.119437 0.219187 0.418687 ;
  RECT 0.200812 0.418687 0.219187 0.437063 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.261188 0.522375 ;
  RECT 0.261188 0.485625 0.300563 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.300563 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0328125 0.066281 0.242812 0.0859685 ;
  RECT 0.242812 0.066281 0.261188 0.0859685 ;
  RECT 0.242812 0.0859685 0.261188 0.138469 ;
      LAYER M1 ;
  RECT 0.0328125 0.066281 0.242812 0.0859685 ;
  RECT 0.242812 0.066281 0.261188 0.0859685 ;
  RECT 0.242812 0.0859685 0.261188 0.138469 ;
  END
END OAI22_X1

MACRO OAI22_X2
  CLASS core ;
  FOREIGN OAI22_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.294 BY 0.504 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.166 0.168 0.177 0.183   ; 
  RECT 0.166 0.183 0.177 0.306   ; 
  RECT 0.166 0.306 0.177 0.324   ; 
  RECT 0.177 0.306 0.264 0.324   ; 
  RECT 0.264 0.183 0.275 0.306   ; 
  RECT 0.264 0.306 0.275 0.324   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.215 0.168 0.226 0.261   ; 
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.117 0.159 0.128 0.319   ; 
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.044 0.159 0.054 0.336   ; 
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.093 0.253 0.103 0.348   ; 
  RECT 0.093 0.348 0.103 0.366   ; 
  RECT 0.103 0.348 0.142 0.366   ; 
  RECT 0.142 0.111 0.152 0.129   ; 
  RECT 0.142 0.129 0.152 0.182   ; 
  RECT 0.142 0.182 0.152 0.253   ; 
  RECT 0.142 0.253 0.152 0.348   ; 
  RECT 0.142 0.348 0.152 0.366   ; 
  RECT 0.152 0.111 0.240 0.129   ; 
  RECT 0.152 0.348 0.240 0.366   ; 
  RECT 0.240 0.111 0.250 0.129   ; 
  RECT 0.240 0.129 0.250 0.182   ; 
  RECT 0.240 0.348 0.250 0.366   ; 
  RECT 0.250 0.348 0.264 0.366   ; 
  RECT 0.264 0.348 0.275 0.366   ; 
  RECT 0.264 0.366 0.275 0.441   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.004 0.486 0.139 0.522   ; 
  RECT 0.139 0.486 0.250 0.522   ; 
  RECT 0.250 0.486 0.275 0.522   ; 
  RECT 0.275 0.486 0.298 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.004 -0.018 0.298 0.018   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.154 0.396 0.240 0.417   ; 
  RECT 0.240 0.396 0.250 0.417   ; 
  RECT 0.240 0.417 0.250 0.457   ; 
  RECT 0.016 0.065 0.264 0.087   ; 
  RECT 0.264 0.065 0.275 0.087   ; 
  RECT 0.264 0.087 0.275 0.138   ; 
  RECT 0.019 0.402 0.139 0.440   ; 
      LAYER M1 ;
  RECT 0.154 0.396 0.240 0.417   ; 
  RECT 0.240 0.396 0.250 0.417   ; 
  RECT 0.240 0.417 0.250 0.457   ; 
  RECT 0.016 0.065 0.264 0.087   ; 
  RECT 0.264 0.065 0.275 0.087   ; 
  RECT 0.264 0.087 0.275 0.138   ; 
  RECT 0.019 0.402 0.139 0.440   ; 
  END
END OAI22_X2

MACRO OR2_X1
  CLASS core ;
  FOREIGN OR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.252 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.063 0.135187 0.336 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.159469 0.0511875 0.420655 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.200812 0.0748125 0.219187 0.42 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.177187 0.522375 ;
  RECT 0.177187 0.485625 0.258562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.258562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0748125 0.0853125 0.093122 0.2205 ;
  RECT 0.0748125 0.2205 0.093122 0.364875 ;
  RECT 0.0748125 0.364875 0.093122 0.38325 ;
  RECT 0.093122 0.364875 0.158812 0.38325 ;
  RECT 0.158812 0.2205 0.177187 0.364875 ;
  RECT 0.158812 0.364875 0.177187 0.38325 ;
      LAYER M1 ;
  RECT 0.0748125 0.0853125 0.093122 0.2205 ;
  RECT 0.0748125 0.2205 0.093122 0.364875 ;
  RECT 0.0748125 0.364875 0.093122 0.38325 ;
  RECT 0.093122 0.364875 0.158812 0.38325 ;
  RECT 0.158812 0.2205 0.177187 0.364875 ;
  RECT 0.158812 0.364875 0.177187 0.38325 ;
  END
END OR2_X1

MACRO OR2_X2
  CLASS core ;
  FOREIGN OR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.252 BY 0.504 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.064 0.159 0.080 0.336   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.028 0.168 0.044 0.336   ; 
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.170 0.042 0.172 0.089   ; 
  RECT 0.170 0.419 0.172 0.462   ; 
  RECT 0.172 0.042 0.188 0.089   ; 
  RECT 0.172 0.089 0.188 0.419   ; 
  RECT 0.172 0.419 0.188 0.462   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.006 0.486 0.152 0.522   ; 
  RECT 0.152 0.486 0.258 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.006 -0.018 0.258 0.018   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.043 0.101 0.082 0.123   ; 
  RECT 0.082 0.101 0.136 0.123   ; 
  RECT 0.082 0.381 0.136 0.399   ; 
  RECT 0.136 0.101 0.152 0.123   ; 
  RECT 0.136 0.123 0.152 0.381   ; 
  RECT 0.136 0.381 0.152 0.399   ; 
      LAYER M1 ;
  RECT 0.043 0.101 0.082 0.123   ; 
  RECT 0.082 0.101 0.136 0.123   ; 
  RECT 0.082 0.381 0.136 0.399   ; 
  RECT 0.136 0.101 0.152 0.123   ; 
  RECT 0.136 0.123 0.152 0.381   ; 
  RECT 0.136 0.381 0.152 0.399   ; 
  END
END OR2_X2

MACRO OR3_X1
  CLASS core ;
  FOREIGN OR3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.336 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.200812 0.126 0.219187 0.378 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.1155 0.126 0.1365 0.378 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0295312 0.126 0.054469 0.378 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.284813 0.0748125 0.303187 0.429187 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.153562 0.522375 ;
  RECT 0.153562 0.485625 0.261188 0.522375 ;
  RECT 0.261188 0.485625 0.342562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.342562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0354375 0.0715315 0.182437 0.089906 ;
  RECT 0.182437 0.0715315 0.242812 0.089906 ;
  RECT 0.182437 0.414095 0.242812 0.441655 ;
  RECT 0.242812 0.0715315 0.261188 0.089906 ;
  RECT 0.242812 0.089906 0.261188 0.414095 ;
  RECT 0.242812 0.414095 0.261188 0.441655 ;
  RECT 0.056372 0.417375 0.153562 0.438375 ;
      LAYER M1 ;
  RECT 0.0354375 0.0715315 0.182437 0.089906 ;
  RECT 0.182437 0.0715315 0.242812 0.089906 ;
  RECT 0.182437 0.414095 0.242812 0.441655 ;
  RECT 0.242812 0.0715315 0.261188 0.089906 ;
  RECT 0.242812 0.089906 0.261188 0.414095 ;
  RECT 0.242812 0.414095 0.261188 0.441655 ;
  RECT 0.056372 0.417375 0.153562 0.438375 ;
  END
END OR3_X1

MACRO OR3_X2
  CLASS core ;
  FOREIGN OR3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.336 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.167344 0.093122 0.294 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.168 0.0511875 0.345187 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.151594 0.177187 0.294 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.240187 0.042 0.242812 0.0853125 ;
  RECT 0.240187 0.417375 0.242812 0.462 ;
  RECT 0.242812 0.042 0.261188 0.0853125 ;
  RECT 0.242812 0.0853125 0.261188 0.417375 ;
  RECT 0.242812 0.417375 0.261188 0.462 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.198187 0.522375 ;
  RECT 0.198187 0.485625 0.219187 0.522375 ;
  RECT 0.219187 0.485625 0.342562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.342562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0328125 0.375965 0.0511875 0.39572 ;
  RECT 0.0328125 0.39572 0.0511875 0.450188 ;
  RECT 0.0511875 0.375965 0.198187 0.39572 ;
  RECT 0.039375 0.101719 0.0924655 0.122719 ;
  RECT 0.0924655 0.101719 0.200812 0.122719 ;
  RECT 0.0924655 0.331405 0.200812 0.352405 ;
  RECT 0.200812 0.101719 0.219187 0.122719 ;
  RECT 0.200812 0.122719 0.219187 0.331405 ;
  RECT 0.200812 0.331405 0.219187 0.352405 ;
      LAYER M1 ;
  RECT 0.0328125 0.375965 0.0511875 0.39572 ;
  RECT 0.0328125 0.39572 0.0511875 0.450188 ;
  RECT 0.0511875 0.375965 0.198187 0.39572 ;
  RECT 0.039375 0.101719 0.0924655 0.122719 ;
  RECT 0.0924655 0.101719 0.200812 0.122719 ;
  RECT 0.0924655 0.331405 0.200812 0.352405 ;
  RECT 0.200812 0.101719 0.219187 0.122719 ;
  RECT 0.200812 0.122719 0.219187 0.331405 ;
  RECT 0.200812 0.331405 0.219187 0.352405 ;
  END
END OR3_X2

MACRO OR4_X1
  CLASS core ;
  FOREIGN OR4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.378 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.242812 0.126 0.261188 0.378 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.1575 0.126 0.1785 0.378 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.129937 0.093122 0.378 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.126 0.0511875 0.378 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.326813 0.0748125 0.345187 0.42 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.195562 0.522375 ;
  RECT 0.195562 0.485625 0.303187 0.522375 ;
  RECT 0.303187 0.485625 0.384562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.384562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0354375 0.066872 0.221812 0.0853125 ;
  RECT 0.221812 0.066872 0.284813 0.0853125 ;
  RECT 0.221812 0.413438 0.284813 0.434437 ;
  RECT 0.284813 0.066872 0.303187 0.0853125 ;
  RECT 0.284813 0.0853125 0.303187 0.413438 ;
  RECT 0.284813 0.413438 0.303187 0.434437 ;
  RECT 0.0958125 0.404905 0.195562 0.429845 ;
      LAYER M1 ;
  RECT 0.0354375 0.066872 0.221812 0.0853125 ;
  RECT 0.221812 0.066872 0.284813 0.0853125 ;
  RECT 0.221812 0.413438 0.284813 0.434437 ;
  RECT 0.284813 0.066872 0.303187 0.0853125 ;
  RECT 0.284813 0.0853125 0.303187 0.413438 ;
  RECT 0.284813 0.413438 0.303187 0.434437 ;
  RECT 0.0958125 0.404905 0.195562 0.429845 ;
  END
END OR4_X1

MACRO OR4_X2
  CLASS core ;
  FOREIGN OR4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.378 BY 0.504 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.181 0.126 0.197 0.348   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.143 0.140 0.159 0.378   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.067 0.140 0.084 0.378   ; 
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.030 0.125 0.046 0.378   ; 
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.293 0.084 0.312 0.462   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.006 0.486 0.178 0.522   ; 
  RECT 0.178 0.486 0.272 0.522   ; 
  RECT 0.272 0.486 0.384 0.522   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.006 -0.018 0.384 0.018   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.086 0.409 0.178 0.447   ; 
  RECT 0.032 0.057 0.202 0.095   ; 
  RECT 0.202 0.057 0.255 0.095   ; 
  RECT 0.202 0.373 0.255 0.409   ; 
  RECT 0.255 0.057 0.272 0.095   ; 
  RECT 0.255 0.095 0.272 0.373   ; 
  RECT 0.255 0.373 0.272 0.409   ; 
      LAYER M1 ;
  RECT 0.086 0.409 0.178 0.447   ; 
  RECT 0.032 0.057 0.202 0.095   ; 
  RECT 0.202 0.057 0.255 0.095   ; 
  RECT 0.202 0.373 0.255 0.409   ; 
  RECT 0.255 0.057 0.272 0.095   ; 
  RECT 0.255 0.095 0.272 0.373   ; 
  RECT 0.255 0.373 0.272 0.409   ; 
  END
END OR4_X2



MACRO TIEH
  CLASS core ;
  FOREIGN TIEH 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.126 BY 0.504 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0715315 0.310405 0.093122 0.462 ;
  RECT 0.093122 0.310405 0.096469 0.462 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.093122 0.522375 ;
  RECT 0.093122 0.485625 0.132562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.132562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0748125 0.063 0.093122 0.28153 ;
      LAYER M1 ;
  RECT 0.0748125 0.063 0.093122 0.28153 ;
  END
END TIEH

MACRO TIEL
  CLASS core ;
  FOREIGN TIEL 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.126 BY 0.504 ;
  PIN Z
    DIRECTION INOUT ;
    PORT
      LAYER M1 ;
  RECT 0.0715315 0.042 0.096469 0.174562 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.093122 0.522375 ;
  RECT 0.093122 0.485625 0.132562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.132562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0748125 0.2205 0.093122 0.441 ;
      LAYER M1 ;
  RECT 0.0748125 0.2205 0.093122 0.441 ;
  END
END TIEL

MACRO XNOR2_X1
  CLASS core ;
  FOREIGN XNOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.378 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.165375 0.137812 0.18375 ;
  RECT 0.116812 0.18375 0.137812 0.280875 ;
  RECT 0.137812 0.165375 0.242812 0.18375 ;
  RECT 0.242812 0.165375 0.261188 0.18375 ;
  RECT 0.242812 0.18375 0.261188 0.280875 ;
  RECT 0.242812 0.280875 0.261188 0.294 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.158812 0.0511875 0.21 ;
  RECT 0.0328125 0.21 0.0511875 0.443625 ;
  RECT 0.0328125 0.443625 0.0511875 0.462 ;
  RECT 0.0511875 0.443625 0.179812 0.462 ;
  RECT 0.179812 0.443625 0.326813 0.462 ;
  RECT 0.326813 0.21 0.345187 0.443625 ;
  RECT 0.326813 0.443625 0.345187 0.462 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.182437 0.358312 0.198187 0.35897 ;
  RECT 0.182437 0.35897 0.198187 0.394405 ;
  RECT 0.182437 0.394405 0.198187 0.395062 ;
  RECT 0.198187 0.108937 0.219187 0.127312 ;
  RECT 0.198187 0.358312 0.219187 0.35897 ;
  RECT 0.198187 0.35897 0.219187 0.394405 ;
  RECT 0.198187 0.394405 0.219187 0.395062 ;
  RECT 0.219187 0.108937 0.284813 0.127312 ;
  RECT 0.219187 0.35897 0.284813 0.394405 ;
  RECT 0.284813 0.108937 0.303187 0.127312 ;
  RECT 0.284813 0.16275 0.303187 0.181125 ;
  RECT 0.284813 0.181125 0.303187 0.358312 ;
  RECT 0.284813 0.358312 0.303187 0.35897 ;
  RECT 0.284813 0.35897 0.303187 0.394405 ;
  RECT 0.303187 0.108937 0.32353 0.127312 ;
  RECT 0.303187 0.16275 0.32353 0.181125 ;
  RECT 0.32353 0.108937 0.34847 0.127312 ;
  RECT 0.32353 0.127312 0.34847 0.16275 ;
  RECT 0.32353 0.16275 0.34847 0.181125 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.179812 0.522375 ;
  RECT 0.179812 0.485625 0.351095 0.522375 ;
  RECT 0.351095 0.485625 0.384562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.384562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.137812 0.066872 0.351095 0.0853125 ;
  RECT 0.0748125 0.12075 0.093122 0.14175 ;
  RECT 0.0748125 0.14175 0.093122 0.223125 ;
  RECT 0.0748125 0.223125 0.093122 0.3045 ;
  RECT 0.0748125 0.3045 0.093122 0.322875 ;
  RECT 0.0748125 0.322875 0.093122 0.36225 ;
  RECT 0.093122 0.12075 0.153562 0.14175 ;
  RECT 0.093122 0.3045 0.153562 0.322875 ;
  RECT 0.153562 0.3045 0.161437 0.322875 ;
  RECT 0.161437 0.223125 0.179812 0.3045 ;
  RECT 0.161437 0.3045 0.179812 0.322875 ;
      LAYER M1 ;
  RECT 0.137812 0.066872 0.351095 0.0853125 ;
  RECT 0.0748125 0.12075 0.093122 0.14175 ;
  RECT 0.0748125 0.14175 0.093122 0.223125 ;
  RECT 0.0748125 0.223125 0.093122 0.3045 ;
  RECT 0.0748125 0.3045 0.093122 0.322875 ;
  RECT 0.0748125 0.322875 0.093122 0.36225 ;
  RECT 0.093122 0.12075 0.153562 0.14175 ;
  RECT 0.093122 0.3045 0.153562 0.322875 ;
  RECT 0.153562 0.3045 0.161437 0.322875 ;
  RECT 0.161437 0.223125 0.179812 0.3045 ;
  RECT 0.161437 0.3045 0.179812 0.322875 ;
  END
END XNOR2_X1

MACRO XOR2_X1
  CLASS core ;
  FOREIGN XOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.378 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.225684 0.137812 0.318937 ;
  RECT 0.116812 0.318937 0.137812 0.337313 ;
  RECT 0.137812 0.318937 0.179812 0.337313 ;
  RECT 0.179812 0.318937 0.242812 0.337313 ;
  RECT 0.242812 0.21 0.261188 0.225684 ;
  RECT 0.242812 0.225684 0.261188 0.318937 ;
  RECT 0.242812 0.318937 0.261188 0.337313 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.042 0.0511875 0.060375 ;
  RECT 0.0328125 0.060375 0.0511875 0.294 ;
  RECT 0.0328125 0.294 0.0511875 0.345187 ;
  RECT 0.0511875 0.042 0.326813 0.060375 ;
  RECT 0.326813 0.042 0.345187 0.060375 ;
  RECT 0.326813 0.060375 0.345187 0.294 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.180469 0.106969 0.206719 0.107625 ;
  RECT 0.180469 0.107625 0.206719 0.145687 ;
  RECT 0.206719 0.106969 0.219187 0.107625 ;
  RECT 0.206719 0.107625 0.219187 0.145687 ;
  RECT 0.206719 0.376688 0.219187 0.395062 ;
  RECT 0.219187 0.107625 0.284813 0.145687 ;
  RECT 0.219187 0.376688 0.284813 0.395062 ;
  RECT 0.284813 0.107625 0.303187 0.145687 ;
  RECT 0.284813 0.145687 0.303187 0.322875 ;
  RECT 0.284813 0.322875 0.303187 0.34125 ;
  RECT 0.284813 0.376688 0.303187 0.395062 ;
  RECT 0.303187 0.322875 0.3255 0.34125 ;
  RECT 0.303187 0.376688 0.3255 0.395062 ;
  RECT 0.3255 0.322875 0.3465 0.34125 ;
  RECT 0.3255 0.34125 0.3465 0.376688 ;
  RECT 0.3255 0.376688 0.3465 0.395062 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.351095 0.522375 ;
  RECT 0.351095 0.485625 0.384562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.384562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.161437 0.418687 0.351095 0.437063 ;
  RECT 0.0748125 0.08925 0.093122 0.18375 ;
  RECT 0.0748125 0.18375 0.093122 0.202125 ;
  RECT 0.0748125 0.202125 0.093122 0.2835 ;
  RECT 0.0748125 0.2835 0.093122 0.36225 ;
  RECT 0.0748125 0.36225 0.093122 0.38325 ;
  RECT 0.093122 0.18375 0.161437 0.202125 ;
  RECT 0.093122 0.36225 0.161437 0.38325 ;
  RECT 0.161437 0.18375 0.162094 0.202125 ;
  RECT 0.161437 0.202125 0.162094 0.2835 ;
  RECT 0.161437 0.36225 0.162094 0.38325 ;
  RECT 0.162094 0.18375 0.179812 0.202125 ;
  RECT 0.162094 0.202125 0.179812 0.2835 ;
      LAYER M1 ;
  RECT 0.161437 0.418687 0.351095 0.437063 ;
  RECT 0.0748125 0.08925 0.093122 0.18375 ;
  RECT 0.0748125 0.18375 0.093122 0.202125 ;
  RECT 0.0748125 0.202125 0.093122 0.2835 ;
  RECT 0.0748125 0.2835 0.093122 0.36225 ;
  RECT 0.0748125 0.36225 0.093122 0.38325 ;
  RECT 0.093122 0.18375 0.161437 0.202125 ;
  RECT 0.093122 0.36225 0.161437 0.38325 ;
  RECT 0.161437 0.18375 0.162094 0.202125 ;
  RECT 0.161437 0.202125 0.162094 0.2835 ;
  RECT 0.161437 0.36225 0.162094 0.38325 ;
  RECT 0.162094 0.18375 0.179812 0.202125 ;
  RECT 0.162094 0.202125 0.179812 0.2835 ;
  END
END XOR2_X1

END LIBRARY
#
# End of file
#
