VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

SITE CORE_TypTyp_0p4_25
  SYMMETRY y ;
  CLASS core ;
SIZE 0.042 BY 0.384 ; 
END CORE_TypTyp_0p4_25


MACRO AND2_X1
  CLASS core ;
  FOREIGN AND2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.2520 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1150 0.1280 0.1370 0.3480 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.0640 0.0530 0.2620 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1990 0.0570 0.2210 0.3200 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.1770 0.3980 ;
        RECT 0.1770 0.3700 0.2590 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.2590 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0730 0.0810 0.0950 0.0950 ;
         RECT 0.0730 0.0950 0.0950 0.2140 ;
         RECT 0.0730 0.2140 0.0950 0.2720 ;
        RECT 0.0930 0.0810 0.1590 0.0950 ;
         RECT 0.1570 0.0810 0.1790 0.0950 ;
         RECT 0.1570 0.0950 0.1790 0.2140 ;
      LAYER M1 ;
         RECT 0.0730 0.0810 0.0950 0.0950 ;
         RECT 0.0730 0.0950 0.0950 0.2140 ;
         RECT 0.0730 0.2140 0.0950 0.2720 ;
        RECT 0.0930 0.0810 0.1590 0.0950 ;
         RECT 0.1570 0.0810 0.1790 0.0950 ;
         RECT 0.1570 0.0950 0.1790 0.2140 ;
  END
END AND2_X1

MACRO AND2_X2
  CLASS core ;
  FOREIGN AND2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.2940 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1150 0.1280 0.1370 0.2560 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.0300 0.1240 0.0540 0.2600 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1885 0.0320 0.2105 0.0650 ;
         RECT 0.1885 0.3190 0.2105 0.3520 ;
         RECT 0.1990 0.0320 0.2210 0.0650 ;
         RECT 0.1990 0.0650 0.2210 0.3190 ;
         RECT 0.1990 0.3190 0.2210 0.3520 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.1770 0.3980 ;
        RECT 0.1770 0.3700 0.3010 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.3010 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0335 0.2870 0.0555 0.3010 ;
        RECT 0.0540 0.0830 0.1590 0.0970 ;
        RECT 0.0540 0.2870 0.1590 0.3010 ;
         RECT 0.1570 0.0830 0.1790 0.0970 ;
         RECT 0.1570 0.0970 0.1790 0.2870 ;
         RECT 0.1570 0.2870 0.1790 0.3010 ;
      LAYER M1 ;
         RECT 0.0335 0.2870 0.0555 0.3010 ;
        RECT 0.0540 0.0830 0.1590 0.0970 ;
        RECT 0.0540 0.2870 0.1590 0.3010 ;
         RECT 0.1570 0.0830 0.1790 0.0970 ;
         RECT 0.1570 0.0970 0.1790 0.2870 ;
         RECT 0.1570 0.2870 0.1790 0.3010 ;
  END
END AND2_X2

MACRO AND3_X1
  CLASS core ;
  FOREIGN AND3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.3360 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1990 0.0960 0.2210 0.2880 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1130 0.0960 0.1380 0.2880 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.0960 0.0530 0.2880 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.2830 0.0570 0.3050 0.3270 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.2610 0.3980 ;
        RECT 0.2610 0.3700 0.3430 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.3430 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.0520 0.0500 0.1560 0.0660 ;
        RECT 0.0350 0.3160 0.1800 0.3300 ;
        RECT 0.1800 0.0480 0.2430 0.0680 ;
        RECT 0.1800 0.3160 0.2430 0.3300 ;
         RECT 0.2410 0.0480 0.2630 0.0680 ;
         RECT 0.2410 0.0680 0.2630 0.3160 ;
         RECT 0.2410 0.3160 0.2630 0.3300 ;
      LAYER M1 ;
        RECT 0.0520 0.0500 0.1560 0.0660 ;
        RECT 0.0350 0.3160 0.1800 0.3300 ;
        RECT 0.1800 0.0480 0.2430 0.0680 ;
        RECT 0.1800 0.3160 0.2430 0.3300 ;
         RECT 0.2410 0.0480 0.2630 0.0680 ;
         RECT 0.2410 0.0680 0.2630 0.3160 ;
         RECT 0.2410 0.3160 0.2630 0.3300 ;
  END
END AND3_X1

MACRO AND3_X2
  CLASS core ;
  FOREIGN AND3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.3360 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1150 0.1600 0.1370 0.2560 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.0300 0.1280 0.0540 0.2560 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1570 0.1510 0.1790 0.2680 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.2305 0.0320 0.2525 0.0780 ;
         RECT 0.2305 0.3190 0.2525 0.3520 ;
         RECT 0.2410 0.0320 0.2630 0.0780 ;
         RECT 0.2410 0.0780 0.2630 0.3190 ;
         RECT 0.2410 0.3190 0.2630 0.3520 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.2190 0.3980 ;
        RECT 0.2190 0.3700 0.3430 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.3430 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0310 0.0360 0.0530 0.0780 ;
         RECT 0.0310 0.0780 0.0530 0.0940 ;
        RECT 0.0520 0.0780 0.1960 0.0940 ;
        RECT 0.0350 0.2900 0.0960 0.3060 ;
        RECT 0.0960 0.1120 0.2010 0.1260 ;
        RECT 0.0960 0.2900 0.2010 0.3060 ;
         RECT 0.1990 0.1120 0.2210 0.1260 ;
         RECT 0.1990 0.1260 0.2210 0.2900 ;
         RECT 0.1990 0.2900 0.2210 0.3060 ;
      LAYER M1 ;
         RECT 0.0310 0.0360 0.0530 0.0780 ;
         RECT 0.0310 0.0780 0.0530 0.0940 ;
        RECT 0.0520 0.0780 0.1960 0.0940 ;
        RECT 0.0350 0.2900 0.0960 0.3060 ;
        RECT 0.0960 0.1120 0.2010 0.1260 ;
        RECT 0.0960 0.2900 0.2010 0.3060 ;
         RECT 0.1990 0.1120 0.2210 0.1260 ;
         RECT 0.1990 0.1260 0.2210 0.2900 ;
         RECT 0.1990 0.2900 0.2210 0.3060 ;
  END
END AND3_X2

MACRO AND4_X1
  CLASS core ;
  FOREIGN AND4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.3780 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.2410 0.0960 0.2630 0.2880 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1575 0.0960 0.1795 0.2880 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.0960 0.0950 0.2560 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.0960 0.0530 0.2880 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.3250 0.0570 0.3470 0.3270 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.3030 0.3980 ;
        RECT 0.3030 0.3700 0.3850 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.3850 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.0540 0.3180 0.2220 0.3340 ;
        RECT 0.2220 0.0500 0.2850 0.0660 ;
        RECT 0.2220 0.3180 0.2850 0.3340 ;
         RECT 0.2830 0.0500 0.3050 0.0660 ;
         RECT 0.2830 0.0660 0.3050 0.3180 ;
         RECT 0.2830 0.3180 0.3050 0.3340 ;
        RECT 0.0920 0.0500 0.1960 0.0740 ;
      LAYER M1 ;
        RECT 0.0540 0.3180 0.2220 0.3340 ;
        RECT 0.2220 0.0500 0.2850 0.0660 ;
        RECT 0.2220 0.3180 0.2850 0.3340 ;
         RECT 0.2830 0.0500 0.3050 0.0660 ;
         RECT 0.2830 0.0660 0.3050 0.3180 ;
         RECT 0.2830 0.3180 0.3050 0.3340 ;
        RECT 0.0920 0.0500 0.1960 0.0740 ;
  END
END AND4_X1

MACRO AND4_X2
  CLASS core ;
  FOREIGN AND4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.4200 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.2410 0.1200 0.2630 0.2880 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1570 0.0960 0.1790 0.2880 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.0960 0.0950 0.2880 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.0960 0.0530 0.2880 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.3250 0.0480 0.3470 0.3200 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.3030 0.3980 ;
        RECT 0.3030 0.3700 0.4270 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.4270 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.0930 0.0500 0.1960 0.0660 ;
        RECT 0.0540 0.3180 0.2240 0.3340 ;
        RECT 0.2240 0.0820 0.2850 0.0980 ;
        RECT 0.2240 0.3180 0.2850 0.3340 ;
         RECT 0.2830 0.0820 0.3050 0.0980 ;
         RECT 0.2830 0.0980 0.3050 0.3180 ;
         RECT 0.2830 0.3180 0.3050 0.3340 ;
      LAYER M1 ;
        RECT 0.0930 0.0500 0.1960 0.0660 ;
        RECT 0.0540 0.3180 0.2240 0.3340 ;
        RECT 0.2240 0.0820 0.2850 0.0980 ;
        RECT 0.2240 0.3180 0.2850 0.3340 ;
         RECT 0.2830 0.0820 0.3050 0.0980 ;
         RECT 0.2830 0.0980 0.3050 0.3180 ;
         RECT 0.2830 0.3180 0.3050 0.3340 ;
  END
END AND4_X2

MACRO ANTENNA
  CLASS core ;
  FOREIGN ANTENNA 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.1260 BY 0.3840 ;
END ANTENNA

MACRO AOI21_X1
  CLASS core ;
  FOREIGN AOI21_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.2520 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1150 0.0960 0.1370 0.2560 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.0670 0.0530 0.2560 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1990 0.0960 0.2210 0.2560 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.0500 0.0950 0.0660 ;
         RECT 0.0730 0.0660 0.0950 0.2680 ;
        RECT 0.0930 0.0500 0.2010 0.0660 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.1960 0.3980 ;
        RECT 0.1960 0.3700 0.2590 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.2590 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0310 0.2900 0.0530 0.3060 ;
         RECT 0.0310 0.3060 0.0530 0.3520 ;
        RECT 0.0520 0.2900 0.1960 0.3060 ;
      LAYER M1 ;
         RECT 0.0310 0.2900 0.0530 0.3060 ;
         RECT 0.0310 0.3060 0.0530 0.3520 ;
        RECT 0.0520 0.2900 0.1960 0.3060 ;
  END
END AOI21_X1

MACRO AOI21_X2
  CLASS core ;
  FOREIGN AOI21_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.3780 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.2410 0.1510 0.2630 0.2240 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1570 0.1150 0.1790 0.1290 ;
         RECT 0.1570 0.1290 0.1790 0.2240 ;
         RECT 0.1570 0.2240 0.1790 0.2560 ;
        RECT 0.1770 0.1150 0.3240 0.1290 ;
        RECT 0.3240 0.1150 0.3480 0.1290 ;
        RECT 0.3240 0.1290 0.3480 0.2240 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.1280 0.0950 0.2240 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.0510 0.0830 0.1170 0.0970 ;
         RECT 0.1150 0.0830 0.1370 0.0970 ;
         RECT 0.1150 0.0970 0.1370 0.2440 ;
         RECT 0.1150 0.2440 0.1370 0.2850 ;
         RECT 0.1150 0.2850 0.1370 0.3000 ;
        RECT 0.1350 0.0830 0.2820 0.0970 ;
        RECT 0.1350 0.2850 0.2820 0.3000 ;
         RECT 0.2725 0.2850 0.2945 0.3000 ;
         RECT 0.2830 0.2440 0.3050 0.2850 ;
         RECT 0.2830 0.2850 0.3050 0.3000 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.3450 0.3980 ;
         RECT 0.3370 0.3700 0.3590 0.3980 ;
        RECT 0.3510 0.3700 0.3850 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.3850 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0310 0.2750 0.0530 0.3180 ;
         RECT 0.0310 0.3180 0.0530 0.3340 ;
        RECT 0.0520 0.3180 0.3270 0.3340 ;
         RECT 0.3250 0.2580 0.3470 0.2750 ;
         RECT 0.3250 0.2750 0.3470 0.3180 ;
         RECT 0.3250 0.3180 0.3470 0.3340 ;
        RECT 0.0960 0.0510 0.3510 0.0650 ;
      LAYER M1 ;
         RECT 0.0310 0.2750 0.0530 0.3180 ;
         RECT 0.0310 0.3180 0.0530 0.3340 ;
        RECT 0.0520 0.3180 0.3270 0.3340 ;
         RECT 0.3250 0.2580 0.3470 0.2750 ;
         RECT 0.3250 0.2750 0.3470 0.3180 ;
         RECT 0.3250 0.3180 0.3470 0.3340 ;
        RECT 0.0960 0.0510 0.3510 0.0650 ;
  END
END AOI21_X2

MACRO AOI22_X1
  CLASS core ;
  FOREIGN AOI22_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.2940 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1570 0.0960 0.1790 0.2560 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.2410 0.0960 0.2630 0.2420 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.0990 0.0950 0.2880 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.0960 0.0530 0.2880 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.0920 0.0510 0.2010 0.0650 ;
         RECT 0.1990 0.0510 0.2210 0.0650 ;
         RECT 0.1990 0.0650 0.2210 0.2910 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.2610 0.3980 ;
        RECT 0.2610 0.3700 0.3010 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.3010 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.0540 0.3150 0.2430 0.3370 ;
         RECT 0.2410 0.2760 0.2630 0.3150 ;
         RECT 0.2410 0.3150 0.2630 0.3370 ;
      LAYER M1 ;
        RECT 0.0540 0.3150 0.2430 0.3370 ;
         RECT 0.2410 0.2760 0.2630 0.3150 ;
         RECT 0.2410 0.3150 0.2630 0.3370 ;
  END
END AOI22_X1

MACRO AOI22_X2
  CLASS core ;
  FOREIGN AOI22_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.5040 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.2830 0.1370 0.3050 0.1510 ;
         RECT 0.2830 0.1510 0.3050 0.2440 ;
         RECT 0.2830 0.2440 0.3050 0.2560 ;
        RECT 0.3030 0.1370 0.4290 0.1510 ;
        RECT 0.4290 0.1370 0.4530 0.1510 ;
         RECT 0.4510 0.1370 0.4730 0.1510 ;
         RECT 0.4510 0.1510 0.4730 0.2440 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.3670 0.1850 0.3890 0.2560 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1990 0.1530 0.2210 0.2630 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1210 0.0530 0.2560 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1570 0.1000 0.1790 0.1140 ;
         RECT 0.1570 0.1140 0.1790 0.1600 ;
        RECT 0.1770 0.1000 0.2380 0.1140 ;
         RECT 0.2295 0.1000 0.2515 0.1140 ;
         RECT 0.2410 0.1000 0.2630 0.1140 ;
         RECT 0.2410 0.1140 0.2630 0.1600 ;
         RECT 0.2410 0.1600 0.2630 0.2320 ;
         RECT 0.2410 0.2320 0.2630 0.2840 ;
         RECT 0.2410 0.2840 0.2630 0.3010 ;
        RECT 0.2610 0.1000 0.4110 0.1140 ;
        RECT 0.2610 0.2840 0.4110 0.3010 ;
         RECT 0.4090 0.1000 0.4310 0.1140 ;
         RECT 0.4090 0.2320 0.4310 0.2840 ;
         RECT 0.4090 0.2840 0.4310 0.3010 ;
        RECT 0.4290 0.1000 0.4530 0.1140 ;
         RECT 0.4510 0.0480 0.4730 0.1000 ;
         RECT 0.4510 0.1000 0.4730 0.1140 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.4710 0.3980 ;
        RECT 0.4710 0.3700 0.5110 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.5110 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.2660 0.0660 0.4110 0.0820 ;
         RECT 0.4090 0.0360 0.4310 0.0660 ;
         RECT 0.4090 0.0660 0.4310 0.0820 ;
        RECT 0.0510 0.3190 0.4530 0.3330 ;
         RECT 0.4510 0.2780 0.4730 0.3190 ;
         RECT 0.4510 0.3190 0.4730 0.3330 ;
        RECT 0.0560 0.0430 0.2380 0.0720 ;
      LAYER M1 ;
        RECT 0.2660 0.0660 0.4110 0.0820 ;
         RECT 0.4090 0.0360 0.4310 0.0660 ;
         RECT 0.4090 0.0660 0.4310 0.0820 ;
        RECT 0.0510 0.3190 0.4530 0.3330 ;
         RECT 0.4510 0.2780 0.4730 0.3190 ;
         RECT 0.4510 0.3190 0.4730 0.3330 ;
        RECT 0.0560 0.0430 0.2380 0.0720 ;
  END
END AOI22_X2

MACRO BUF_X1
  CLASS core ;
  FOREIGN BUF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.2100 BY 0.3840 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.0960 0.0530 0.2880 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1575 0.0570 0.1795 0.3520 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.0940 0.3980 ;
        RECT 0.0940 0.3700 0.2170 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.2170 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0730 0.0360 0.0950 0.0920 ;
         RECT 0.0730 0.0920 0.0950 0.1060 ;
         RECT 0.0730 0.1060 0.0950 0.2140 ;
         RECT 0.0730 0.2140 0.0950 0.2280 ;
         RECT 0.0730 0.2280 0.0950 0.2790 ;
         RECT 0.0825 0.0920 0.1045 0.1060 ;
         RECT 0.0825 0.1060 0.1045 0.2140 ;
         RECT 0.0825 0.2140 0.1045 0.2280 ;
      LAYER M1 ;
         RECT 0.0730 0.0360 0.0950 0.0920 ;
         RECT 0.0730 0.0920 0.0950 0.1060 ;
         RECT 0.0730 0.1060 0.0950 0.2140 ;
         RECT 0.0730 0.2140 0.0950 0.2280 ;
         RECT 0.0730 0.2280 0.0950 0.2790 ;
         RECT 0.0825 0.0920 0.1045 0.1060 ;
         RECT 0.0825 0.1060 0.1045 0.2140 ;
         RECT 0.0825 0.2140 0.1045 0.2280 ;
  END
END BUF_X1

MACRO BUF_X2
  CLASS core ;
  FOREIGN BUF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.2100 BY 0.3840 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1340 0.0530 0.2560 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1040 0.3020 0.1260 0.3520 ;
         RECT 0.1055 0.0360 0.1275 0.0660 ;
         RECT 0.1055 0.3020 0.1275 0.3520 ;
         RECT 0.1150 0.0360 0.1370 0.0660 ;
         RECT 0.1150 0.0660 0.1370 0.3020 ;
         RECT 0.1150 0.3020 0.1370 0.3520 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.0930 0.3980 ;
        RECT 0.0930 0.3700 0.2170 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.2170 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0195 0.2780 0.0415 0.2920 ;
         RECT 0.0195 0.2920 0.0415 0.3430 ;
         RECT 0.0310 0.0480 0.0530 0.0960 ;
         RECT 0.0310 0.0960 0.0530 0.1100 ;
         RECT 0.0310 0.2780 0.0530 0.2920 ;
         RECT 0.0310 0.2920 0.0530 0.3430 ;
         RECT 0.0425 0.0960 0.0645 0.1100 ;
         RECT 0.0425 0.2780 0.0645 0.2920 ;
         RECT 0.0425 0.2920 0.0645 0.3430 ;
         RECT 0.0545 0.0960 0.0765 0.1100 ;
         RECT 0.0545 0.2780 0.0765 0.2920 ;
         RECT 0.0730 0.0960 0.0950 0.1100 ;
         RECT 0.0730 0.1100 0.0950 0.2780 ;
         RECT 0.0730 0.2780 0.0950 0.2920 ;
      LAYER M1 ;
         RECT 0.0195 0.2780 0.0415 0.2920 ;
         RECT 0.0195 0.2920 0.0415 0.3430 ;
         RECT 0.0310 0.0480 0.0530 0.0960 ;
         RECT 0.0310 0.0960 0.0530 0.1100 ;
         RECT 0.0310 0.2780 0.0530 0.2920 ;
         RECT 0.0310 0.2920 0.0530 0.3430 ;
         RECT 0.0425 0.0960 0.0645 0.1100 ;
         RECT 0.0425 0.2780 0.0645 0.2920 ;
         RECT 0.0425 0.2920 0.0645 0.3430 ;
         RECT 0.0545 0.0960 0.0765 0.1100 ;
         RECT 0.0545 0.2780 0.0765 0.2920 ;
         RECT 0.0730 0.0960 0.0950 0.1100 ;
         RECT 0.0730 0.1100 0.0950 0.2780 ;
         RECT 0.0730 0.2780 0.0950 0.2920 ;
  END
END BUF_X2

MACRO BUF_X4
  CLASS core ;
  FOREIGN BUF_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.3360 BY 0.3840 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1150 0.1210 0.1370 0.2630 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.0950 0.0510 0.1380 0.0650 ;
        RECT 0.1380 0.0510 0.1770 0.0650 ;
        RECT 0.1380 0.3190 0.1770 0.3330 ;
        RECT 0.1770 0.0510 0.2420 0.0650 ;
        RECT 0.1770 0.3190 0.2420 0.3330 ;
         RECT 0.2410 0.0510 0.2630 0.0650 ;
         RECT 0.2410 0.0650 0.2630 0.3190 ;
         RECT 0.2410 0.3190 0.2630 0.3330 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.1770 0.3980 ;
        RECT 0.1770 0.3700 0.3430 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.3430 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.0180 0.0830 0.0560 0.0990 ;
        RECT 0.0560 0.0830 0.1590 0.0990 ;
        RECT 0.0560 0.2850 0.1590 0.3010 ;
         RECT 0.1570 0.0830 0.1790 0.0990 ;
         RECT 0.1570 0.0990 0.1790 0.2850 ;
         RECT 0.1570 0.2850 0.1790 0.3010 ;
      LAYER M1 ;
        RECT 0.0180 0.0830 0.0560 0.0990 ;
        RECT 0.0560 0.0830 0.1590 0.0990 ;
        RECT 0.0560 0.2850 0.1590 0.3010 ;
         RECT 0.1570 0.0830 0.1790 0.0990 ;
         RECT 0.1570 0.0990 0.1790 0.2850 ;
         RECT 0.1570 0.2850 0.1790 0.3010 ;
  END
END BUF_X4

MACRO BUF_X8
  CLASS core ;
  FOREIGN BUF_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.5880 BY 0.3840 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1280 0.0530 0.1830 ;
         RECT 0.0310 0.1830 0.0530 0.1990 ;
         RECT 0.0310 0.1990 0.0530 0.2560 ;
        RECT 0.0510 0.1830 0.1960 0.1990 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.2220 0.0510 0.4590 0.0650 ;
        RECT 0.2220 0.3190 0.4590 0.3330 ;
        RECT 0.4590 0.0510 0.4950 0.0650 ;
        RECT 0.4590 0.3190 0.4950 0.3330 ;
         RECT 0.4930 0.0510 0.5150 0.0650 ;
         RECT 0.4930 0.0650 0.5150 0.3190 ;
         RECT 0.4930 0.3190 0.5150 0.3330 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.4590 0.3980 ;
        RECT 0.4590 0.3700 0.5950 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.5950 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0590 0.0490 0.0810 0.0930 ;
         RECT 0.0590 0.0930 0.0810 0.1070 ;
         RECT 0.0730 0.0490 0.0950 0.0930 ;
         RECT 0.0730 0.0930 0.0950 0.1070 ;
         RECT 0.0730 0.2640 0.0950 0.2920 ;
         RECT 0.0730 0.2920 0.0950 0.3350 ;
         RECT 0.0870 0.0490 0.1090 0.0930 ;
         RECT 0.0870 0.0930 0.1090 0.1070 ;
         RECT 0.0870 0.2640 0.1090 0.2920 ;
        RECT 0.1030 0.0930 0.2320 0.1070 ;
        RECT 0.1030 0.2640 0.2320 0.2920 ;
         RECT 0.2305 0.0930 0.2525 0.1070 ;
         RECT 0.2305 0.1070 0.2525 0.1700 ;
         RECT 0.2305 0.1700 0.2525 0.1840 ;
         RECT 0.2305 0.1840 0.2525 0.2640 ;
         RECT 0.2305 0.2640 0.2525 0.2920 ;
        RECT 0.2510 0.1700 0.4590 0.1840 ;
      LAYER M1 ;
         RECT 0.0590 0.0490 0.0810 0.0930 ;
         RECT 0.0590 0.0930 0.0810 0.1070 ;
         RECT 0.0730 0.0490 0.0950 0.0930 ;
         RECT 0.0730 0.0930 0.0950 0.1070 ;
         RECT 0.0730 0.2640 0.0950 0.2920 ;
         RECT 0.0730 0.2920 0.0950 0.3350 ;
         RECT 0.0870 0.0490 0.1090 0.0930 ;
         RECT 0.0870 0.0930 0.1090 0.1070 ;
         RECT 0.0870 0.2640 0.1090 0.2920 ;
        RECT 0.1030 0.0930 0.2320 0.1070 ;
        RECT 0.1030 0.2640 0.2320 0.2920 ;
         RECT 0.2305 0.0930 0.2525 0.1070 ;
         RECT 0.2305 0.1070 0.2525 0.1700 ;
         RECT 0.2305 0.1700 0.2525 0.1840 ;
         RECT 0.2305 0.1840 0.2525 0.2640 ;
         RECT 0.2305 0.2640 0.2525 0.2920 ;
        RECT 0.2510 0.1700 0.4590 0.1840 ;
  END
END BUF_X8

MACRO BUF_X12
  CLASS core ;
  FOREIGN BUF_X12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.8400 BY 0.3840 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1180 0.0530 0.1830 ;
         RECT 0.0310 0.1830 0.0530 0.1990 ;
         RECT 0.0310 0.1990 0.0530 0.2580 ;
        RECT 0.0520 0.1830 0.2800 0.1990 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.3060 0.0510 0.7020 0.0650 ;
        RECT 0.3060 0.3190 0.7020 0.3330 ;
        RECT 0.7020 0.0510 0.7450 0.0650 ;
        RECT 0.7020 0.3190 0.7450 0.3330 ;
         RECT 0.7445 0.0510 0.7665 0.0650 ;
         RECT 0.7445 0.0650 0.7665 0.3190 ;
         RECT 0.7445 0.3190 0.7665 0.3330 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.7020 0.3980 ;
        RECT 0.7020 0.3700 0.8470 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.8470 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0580 0.2760 0.0800 0.2920 ;
         RECT 0.0580 0.2920 0.0800 0.3350 ;
         RECT 0.0730 0.0490 0.0950 0.0920 ;
         RECT 0.0730 0.0920 0.0950 0.1080 ;
         RECT 0.0730 0.2760 0.0950 0.2920 ;
         RECT 0.0730 0.2920 0.0950 0.3350 ;
         RECT 0.0875 0.0920 0.1095 0.1080 ;
         RECT 0.0875 0.2760 0.1095 0.2920 ;
         RECT 0.0875 0.2920 0.1095 0.3350 ;
        RECT 0.1030 0.0920 0.3030 0.1080 ;
        RECT 0.1030 0.2760 0.3030 0.2920 ;
         RECT 0.3015 0.0920 0.3235 0.1080 ;
         RECT 0.3015 0.1080 0.3235 0.1850 ;
         RECT 0.3015 0.1850 0.3235 0.1990 ;
         RECT 0.3015 0.1990 0.3235 0.2760 ;
         RECT 0.3015 0.2760 0.3235 0.2920 ;
        RECT 0.3220 0.1850 0.7020 0.1990 ;
      LAYER M1 ;
         RECT 0.0580 0.2760 0.0800 0.2920 ;
         RECT 0.0580 0.2920 0.0800 0.3350 ;
         RECT 0.0730 0.0490 0.0950 0.0920 ;
         RECT 0.0730 0.0920 0.0950 0.1080 ;
         RECT 0.0730 0.2760 0.0950 0.2920 ;
         RECT 0.0730 0.2920 0.0950 0.3350 ;
         RECT 0.0875 0.0920 0.1095 0.1080 ;
         RECT 0.0875 0.2760 0.1095 0.2920 ;
         RECT 0.0875 0.2920 0.1095 0.3350 ;
        RECT 0.1030 0.0920 0.3030 0.1080 ;
        RECT 0.1030 0.2760 0.3030 0.2920 ;
         RECT 0.3015 0.0920 0.3235 0.1080 ;
         RECT 0.3015 0.1080 0.3235 0.1850 ;
         RECT 0.3015 0.1850 0.3235 0.1990 ;
         RECT 0.3015 0.1990 0.3235 0.2760 ;
         RECT 0.3015 0.2760 0.3235 0.2920 ;
        RECT 0.3220 0.1850 0.7020 0.1990 ;
  END
END BUF_X12

MACRO BUF_X16
  CLASS core ;
  FOREIGN BUF_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 1.0920 BY 0.3840 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1160 0.0530 0.1780 ;
         RECT 0.0310 0.1780 0.0530 0.2060 ;
         RECT 0.0310 0.2060 0.0530 0.2560 ;
        RECT 0.0510 0.1780 0.3640 0.2060 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.3900 0.0510 0.9540 0.0650 ;
        RECT 0.3900 0.3160 0.9540 0.3300 ;
        RECT 0.9540 0.0510 0.9980 0.0650 ;
        RECT 0.9540 0.3160 0.9980 0.3300 ;
         RECT 0.9970 0.0510 1.0190 0.0650 ;
         RECT 0.9970 0.0650 1.0190 0.3160 ;
         RECT 0.9970 0.3160 1.0190 0.3300 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.9540 0.3980 ;
        RECT 0.9540 0.3700 1.0990 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 1.0990 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0730 0.0490 0.0950 0.1020 ;
         RECT 0.0730 0.1020 0.0950 0.1160 ;
         RECT 0.0730 0.2290 0.0950 0.2430 ;
         RECT 0.0730 0.2430 0.0950 0.3220 ;
        RECT 0.0930 0.1020 0.3870 0.1160 ;
        RECT 0.0930 0.2290 0.3870 0.2430 ;
         RECT 0.3855 0.1020 0.4075 0.1160 ;
         RECT 0.3855 0.1160 0.4075 0.1840 ;
         RECT 0.3855 0.1840 0.4075 0.1980 ;
         RECT 0.3855 0.1980 0.4075 0.2290 ;
         RECT 0.3855 0.2290 0.4075 0.2430 ;
        RECT 0.4060 0.1840 0.9540 0.1980 ;
      LAYER M1 ;
         RECT 0.0730 0.0490 0.0950 0.1020 ;
         RECT 0.0730 0.1020 0.0950 0.1160 ;
         RECT 0.0730 0.2290 0.0950 0.2430 ;
         RECT 0.0730 0.2430 0.0950 0.3220 ;
        RECT 0.0930 0.1020 0.3870 0.1160 ;
        RECT 0.0930 0.2290 0.3870 0.2430 ;
         RECT 0.3855 0.1020 0.4075 0.1160 ;
         RECT 0.3855 0.1160 0.4075 0.1840 ;
         RECT 0.3855 0.1840 0.4075 0.1980 ;
         RECT 0.3855 0.1980 0.4075 0.2290 ;
         RECT 0.3855 0.2290 0.4075 0.2430 ;
        RECT 0.4060 0.1840 0.9540 0.1980 ;
  END
END BUF_X16

MACRO CLKBUF_X1
  CLASS core ;
  FOREIGN CLKBUF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.2100 BY 0.3840 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.0960 0.0530 0.2880 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1575 0.0570 0.1795 0.3520 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.0940 0.3980 ;
        RECT 0.0940 0.3700 0.2170 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.2170 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0730 0.0360 0.0950 0.0920 ;
         RECT 0.0730 0.0920 0.0950 0.1060 ;
         RECT 0.0730 0.1060 0.0950 0.1960 ;
         RECT 0.0730 0.1960 0.0950 0.2290 ;
         RECT 0.0730 0.2290 0.0950 0.2620 ;
         RECT 0.0825 0.0920 0.1045 0.1060 ;
         RECT 0.0825 0.1060 0.1045 0.1960 ;
         RECT 0.0825 0.1960 0.1045 0.2290 ;
      LAYER M1 ;
         RECT 0.0730 0.0360 0.0950 0.0920 ;
         RECT 0.0730 0.0920 0.0950 0.1060 ;
         RECT 0.0730 0.1060 0.0950 0.1960 ;
         RECT 0.0730 0.1960 0.0950 0.2290 ;
         RECT 0.0730 0.2290 0.0950 0.2620 ;
         RECT 0.0825 0.0920 0.1045 0.1060 ;
         RECT 0.0825 0.1060 0.1045 0.1960 ;
         RECT 0.0825 0.1960 0.1045 0.2290 ;
  END
END CLKBUF_X1

MACRO CLKBUF_X2
  CLASS core ;
  FOREIGN CLKBUF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.2100 BY 0.3840 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1480 0.0530 0.2560 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1045 0.3190 0.1265 0.3520 ;
         RECT 0.1150 0.0360 0.1370 0.3190 ;
         RECT 0.1150 0.3190 0.1370 0.3520 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.0930 0.3980 ;
        RECT 0.0930 0.3700 0.2170 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.2170 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0310 0.0640 0.0530 0.0960 ;
         RECT 0.0310 0.0960 0.0530 0.1100 ;
         RECT 0.0310 0.2780 0.0530 0.2920 ;
         RECT 0.0310 0.2920 0.0530 0.3430 ;
        RECT 0.0520 0.0960 0.0750 0.1100 ;
        RECT 0.0520 0.2780 0.0750 0.2920 ;
         RECT 0.0730 0.0960 0.0950 0.1100 ;
         RECT 0.0730 0.1100 0.0950 0.2780 ;
         RECT 0.0730 0.2780 0.0950 0.2920 ;
      LAYER M1 ;
         RECT 0.0310 0.0640 0.0530 0.0960 ;
         RECT 0.0310 0.0960 0.0530 0.1100 ;
         RECT 0.0310 0.2780 0.0530 0.2920 ;
         RECT 0.0310 0.2920 0.0530 0.3430 ;
        RECT 0.0520 0.0960 0.0750 0.1100 ;
        RECT 0.0520 0.2780 0.0750 0.2920 ;
         RECT 0.0730 0.0960 0.0950 0.1100 ;
         RECT 0.0730 0.1100 0.0950 0.2780 ;
         RECT 0.0730 0.2780 0.0950 0.2920 ;
  END
END CLKBUF_X2

MACRO CLKBUF_X4
  CLASS core ;
  FOREIGN CLKBUF_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.3360 BY 0.3840 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.1210 0.0950 0.2630 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.0950 0.0510 0.1350 0.0650 ;
        RECT 0.1350 0.0510 0.2420 0.0650 ;
        RECT 0.1350 0.3190 0.2420 0.3330 ;
         RECT 0.2410 0.0510 0.2630 0.0650 ;
         RECT 0.2410 0.0650 0.2630 0.3190 ;
         RECT 0.2410 0.3190 0.2630 0.3330 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.1350 0.3980 ;
        RECT 0.1350 0.3700 0.3430 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.3430 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.0270 0.0830 0.0540 0.0970 ;
        RECT 0.0540 0.0830 0.1170 0.0970 ;
        RECT 0.0540 0.2870 0.1170 0.3010 ;
         RECT 0.1150 0.0830 0.1370 0.0970 ;
         RECT 0.1150 0.0970 0.1370 0.2870 ;
         RECT 0.1150 0.2870 0.1370 0.3010 ;
      LAYER M1 ;
        RECT 0.0270 0.0830 0.0540 0.0970 ;
        RECT 0.0540 0.0830 0.1170 0.0970 ;
        RECT 0.0540 0.2870 0.1170 0.3010 ;
         RECT 0.1150 0.0830 0.1370 0.0970 ;
         RECT 0.1150 0.0970 0.1370 0.2870 ;
         RECT 0.1150 0.2870 0.1370 0.3010 ;
  END
END CLKBUF_X4

MACRO CLKBUF_X8
  CLASS core ;
  FOREIGN CLKBUF_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.5880 BY 0.3840 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1280 0.0530 0.1640 ;
         RECT 0.0310 0.1640 0.0530 0.1780 ;
         RECT 0.0310 0.1780 0.0530 0.2560 ;
         RECT 0.0405 0.1280 0.0625 0.1640 ;
         RECT 0.0405 0.1640 0.0625 0.1780 ;
        RECT 0.0520 0.1640 0.2090 0.1780 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.2220 0.0510 0.4710 0.0650 ;
        RECT 0.2220 0.3190 0.4710 0.3330 ;
        RECT 0.4710 0.0510 0.4950 0.0650 ;
        RECT 0.4710 0.3190 0.4950 0.3330 ;
         RECT 0.4930 0.0510 0.5150 0.0650 ;
         RECT 0.4930 0.0650 0.5150 0.3190 ;
         RECT 0.4930 0.3190 0.5150 0.3330 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.4710 0.3980 ;
        RECT 0.4710 0.3700 0.5950 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.5950 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.0330 0.0830 0.0750 0.0970 ;
         RECT 0.0730 0.0830 0.0950 0.0970 ;
         RECT 0.0730 0.2250 0.0950 0.2410 ;
         RECT 0.0730 0.2410 0.0950 0.2710 ;
        RECT 0.0930 0.0830 0.2660 0.0970 ;
        RECT 0.0930 0.2250 0.2660 0.2410 ;
         RECT 0.2645 0.0830 0.2865 0.0970 ;
         RECT 0.2645 0.0970 0.2865 0.1780 ;
         RECT 0.2645 0.1780 0.2865 0.2070 ;
         RECT 0.2645 0.2070 0.2865 0.2250 ;
         RECT 0.2645 0.2250 0.2865 0.2410 ;
        RECT 0.2850 0.1780 0.4710 0.2070 ;
      LAYER M1 ;
        RECT 0.0330 0.0830 0.0750 0.0970 ;
         RECT 0.0730 0.0830 0.0950 0.0970 ;
         RECT 0.0730 0.2250 0.0950 0.2410 ;
         RECT 0.0730 0.2410 0.0950 0.2710 ;
        RECT 0.0930 0.0830 0.2660 0.0970 ;
        RECT 0.0930 0.2250 0.2660 0.2410 ;
         RECT 0.2645 0.0830 0.2865 0.0970 ;
         RECT 0.2645 0.0970 0.2865 0.1780 ;
         RECT 0.2645 0.1780 0.2865 0.2070 ;
         RECT 0.2645 0.2070 0.2865 0.2250 ;
         RECT 0.2645 0.2250 0.2865 0.2410 ;
        RECT 0.2850 0.1780 0.4710 0.2070 ;
  END
END CLKBUF_X8

MACRO CLKBUF_X12
  CLASS core ;
  FOREIGN CLKBUF_X12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.8400 BY 0.3840 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.0300 0.1190 0.0540 0.1680 ;
        RECT 0.0300 0.1680 0.0540 0.1840 ;
        RECT 0.0300 0.1840 0.0540 0.2650 ;
        RECT 0.0540 0.1680 0.2800 0.1840 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.3060 0.0510 0.6550 0.0650 ;
        RECT 0.3060 0.3190 0.6550 0.3330 ;
        RECT 0.6550 0.0510 0.7450 0.0650 ;
        RECT 0.6550 0.3190 0.7450 0.3330 ;
         RECT 0.7445 0.0510 0.7665 0.0650 ;
         RECT 0.7445 0.0650 0.7665 0.3190 ;
         RECT 0.7445 0.3190 0.7665 0.3330 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.6550 0.3980 ;
        RECT 0.6550 0.3700 0.8470 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.8470 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.0280 0.0830 0.0750 0.0970 ;
         RECT 0.0730 0.0830 0.0950 0.0970 ;
         RECT 0.0730 0.2750 0.0950 0.2890 ;
         RECT 0.0730 0.2890 0.0950 0.3350 ;
        RECT 0.0930 0.0830 0.3030 0.0970 ;
        RECT 0.0930 0.2750 0.3030 0.2890 ;
         RECT 0.3015 0.0830 0.3235 0.0970 ;
         RECT 0.3015 0.0970 0.3235 0.1570 ;
         RECT 0.3015 0.1570 0.3235 0.1730 ;
         RECT 0.3015 0.1730 0.3235 0.2750 ;
         RECT 0.3015 0.2750 0.3235 0.2890 ;
         RECT 0.3120 0.0830 0.3340 0.0970 ;
         RECT 0.3120 0.0970 0.3340 0.1570 ;
         RECT 0.3120 0.1570 0.3340 0.1730 ;
        RECT 0.3240 0.1570 0.6550 0.1730 ;
      LAYER M1 ;
        RECT 0.0280 0.0830 0.0750 0.0970 ;
         RECT 0.0730 0.0830 0.0950 0.0970 ;
         RECT 0.0730 0.2750 0.0950 0.2890 ;
         RECT 0.0730 0.2890 0.0950 0.3350 ;
        RECT 0.0930 0.0830 0.3030 0.0970 ;
        RECT 0.0930 0.2750 0.3030 0.2890 ;
         RECT 0.3015 0.0830 0.3235 0.0970 ;
         RECT 0.3015 0.0970 0.3235 0.1570 ;
         RECT 0.3015 0.1570 0.3235 0.1730 ;
         RECT 0.3015 0.1730 0.3235 0.2750 ;
         RECT 0.3015 0.2750 0.3235 0.2890 ;
         RECT 0.3120 0.0830 0.3340 0.0970 ;
         RECT 0.3120 0.0970 0.3340 0.1570 ;
         RECT 0.3120 0.1570 0.3340 0.1730 ;
        RECT 0.3240 0.1570 0.6550 0.1730 ;
  END
END CLKBUF_X12

MACRO CLKBUF_X16
  CLASS core ;
  FOREIGN CLKBUF_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 1.0920 BY 0.3840 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1110 0.0530 0.1630 ;
         RECT 0.0310 0.1630 0.0530 0.1790 ;
         RECT 0.0310 0.1790 0.0530 0.2630 ;
        RECT 0.0510 0.1630 0.3640 0.1790 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.3900 0.0430 0.9540 0.0720 ;
        RECT 0.3900 0.3120 0.9540 0.3400 ;
        RECT 0.9540 0.0430 0.9980 0.0720 ;
        RECT 0.9540 0.3120 0.9980 0.3400 ;
         RECT 0.9970 0.0430 1.0190 0.0720 ;
         RECT 0.9970 0.0720 1.0190 0.3120 ;
         RECT 0.9970 0.3120 1.0190 0.3400 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.9540 0.3980 ;
        RECT 0.9540 0.3700 1.0990 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 1.0990 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0730 0.0540 0.0950 0.1020 ;
         RECT 0.0730 0.1020 0.0950 0.1160 ;
         RECT 0.0730 0.2620 0.0950 0.2810 ;
         RECT 0.0730 0.2810 0.0950 0.3190 ;
        RECT 0.0930 0.1020 0.3900 0.1160 ;
        RECT 0.0930 0.2620 0.3900 0.2810 ;
        RECT 0.3900 0.1020 0.4290 0.1160 ;
        RECT 0.3900 0.1160 0.4290 0.1580 ;
        RECT 0.3900 0.1580 0.4290 0.1720 ;
        RECT 0.3900 0.1720 0.4290 0.2620 ;
        RECT 0.3900 0.2620 0.4290 0.2810 ;
        RECT 0.4290 0.1580 0.9540 0.1720 ;
      LAYER M1 ;
         RECT 0.0730 0.0540 0.0950 0.1020 ;
         RECT 0.0730 0.1020 0.0950 0.1160 ;
         RECT 0.0730 0.2620 0.0950 0.2810 ;
         RECT 0.0730 0.2810 0.0950 0.3190 ;
        RECT 0.0930 0.1020 0.3900 0.1160 ;
        RECT 0.0930 0.2620 0.3900 0.2810 ;
        RECT 0.3900 0.1020 0.4290 0.1160 ;
        RECT 0.3900 0.1160 0.4290 0.1580 ;
        RECT 0.3900 0.1580 0.4290 0.1720 ;
        RECT 0.3900 0.1720 0.4290 0.2620 ;
        RECT 0.3900 0.2620 0.4290 0.2810 ;
        RECT 0.4290 0.1580 0.9540 0.1720 ;
  END
END CLKBUF_X16

MACRO CLKGATETST_X1
  CLASS core ;
  FOREIGN CLKGATETST_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.7140 BY 0.3840 ;
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
         RECT 0.4510 0.1190 0.4730 0.2560 ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.1280 0.0950 0.3360 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1600 0.0530 0.3360 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.6610 0.0480 0.6830 0.3270 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.2400 0.3980 ;
        RECT 0.2400 0.3700 0.5970 0.3980 ;
        RECT 0.5970 0.3700 0.6390 0.3980 ;
        RECT 0.6390 0.3700 0.7210 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.7210 0.0140 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
         RECT 0.1380 0.1960 0.4500 0.2200 ;
         RECT 0.0960 0.2280 0.3430 0.2520 ;
         RECT 0.4790 0.1960 0.6600 0.2200 ;
      LAYER MINT1 ;
         RECT 0.1380 0.1960 0.4500 0.2200 ;
         RECT 0.0960 0.2280 0.3430 0.2520 ;
         RECT 0.4790 0.1960 0.6600 0.2200 ;
      LAYER M1 ;
         RECT 0.0310 0.0510 0.0530 0.0650 ;
         RECT 0.0310 0.0650 0.0530 0.1060 ;
        RECT 0.0520 0.0510 0.1560 0.0650 ;
         RECT 0.1570 0.1320 0.1790 0.2700 ;
         RECT 0.2410 0.1210 0.2630 0.2510 ;
         RECT 0.3025 0.1860 0.3245 0.2550 ;
         RECT 0.4090 0.0830 0.4310 0.0970 ;
         RECT 0.4090 0.0970 0.4310 0.2780 ;
         RECT 0.4090 0.2780 0.4310 0.2960 ;
        RECT 0.4290 0.0830 0.4920 0.0970 ;
        RECT 0.4290 0.2780 0.4920 0.2960 ;
         RECT 0.4825 0.0830 0.5045 0.0970 ;
        RECT 0.4950 0.1240 0.5180 0.2320 ;
        RECT 0.4950 0.2320 0.5180 0.2510 ;
         RECT 0.5165 0.2320 0.5385 0.2510 ;
         RECT 0.5350 0.2320 0.5570 0.2510 ;
         RECT 0.5350 0.2510 0.5570 0.2920 ;
         RECT 0.6190 0.1130 0.6410 0.2870 ;
         RECT 0.1150 0.0830 0.1370 0.0970 ;
         RECT 0.1150 0.0970 0.1370 0.3140 ;
         RECT 0.1150 0.3140 0.1370 0.3380 ;
        RECT 0.1350 0.0830 0.1980 0.0970 ;
        RECT 0.1350 0.3140 0.1980 0.3380 ;
        RECT 0.1980 0.3140 0.2400 0.3380 ;
         RECT 0.1990 0.1540 0.2210 0.2730 ;
         RECT 0.1990 0.2730 0.2210 0.2870 ;
        RECT 0.2190 0.2730 0.3660 0.2870 ;
         RECT 0.3655 0.0920 0.3875 0.1540 ;
         RECT 0.3655 0.1540 0.3875 0.2730 ;
         RECT 0.3655 0.2730 0.3875 0.2870 ;
         RECT 0.2830 0.0510 0.3050 0.0650 ;
         RECT 0.2830 0.0650 0.3050 0.1670 ;
         RECT 0.2935 0.0510 0.3155 0.0650 ;
        RECT 0.3060 0.0510 0.5790 0.0650 ;
        RECT 0.3060 0.3140 0.5790 0.3380 ;
         RECT 0.5770 0.0510 0.5990 0.0650 ;
         RECT 0.5770 0.0650 0.5990 0.1670 ;
         RECT 0.5770 0.1670 0.5990 0.3140 ;
         RECT 0.5770 0.3140 0.5990 0.3380 ;
      LAYER V1 ;
        RECT 0.1170 0.2330 0.1350 0.2470 ;
        RECT 0.1590 0.2010 0.1770 0.2150 ;
        RECT 0.2430 0.2010 0.2610 0.2150 ;
        RECT 0.3030 0.2330 0.3220 0.2470 ;
        RECT 0.4110 0.2010 0.4290 0.2150 ;
        RECT 0.5000 0.2010 0.5180 0.2150 ;
        RECT 0.6210 0.2010 0.6390 0.2150 ;
      LAYER M1 ;
         RECT 0.0310 0.0510 0.0530 0.0650 ;
         RECT 0.0310 0.0650 0.0530 0.1060 ;
        RECT 0.0520 0.0510 0.1560 0.0650 ;
         RECT 0.1570 0.1320 0.1790 0.2700 ;
         RECT 0.2410 0.1210 0.2630 0.2510 ;
         RECT 0.3025 0.1860 0.3245 0.2550 ;
         RECT 0.4090 0.0830 0.4310 0.0970 ;
         RECT 0.4090 0.0970 0.4310 0.2780 ;
         RECT 0.4090 0.2780 0.4310 0.2960 ;
        RECT 0.4290 0.0830 0.4920 0.0970 ;
        RECT 0.4290 0.2780 0.4920 0.2960 ;
         RECT 0.4825 0.0830 0.5045 0.0970 ;
        RECT 0.4950 0.1240 0.5180 0.2320 ;
        RECT 0.4950 0.2320 0.5180 0.2510 ;
         RECT 0.5165 0.2320 0.5385 0.2510 ;
         RECT 0.5350 0.2320 0.5570 0.2510 ;
         RECT 0.5350 0.2510 0.5570 0.2920 ;
         RECT 0.6190 0.1130 0.6410 0.2870 ;
         RECT 0.1150 0.0830 0.1370 0.0970 ;
         RECT 0.1150 0.0970 0.1370 0.3140 ;
         RECT 0.1150 0.3140 0.1370 0.3380 ;
        RECT 0.1350 0.0830 0.1980 0.0970 ;
        RECT 0.1350 0.3140 0.1980 0.3380 ;
        RECT 0.1980 0.3140 0.2400 0.3380 ;
         RECT 0.1990 0.1540 0.2210 0.2730 ;
         RECT 0.1990 0.2730 0.2210 0.2870 ;
        RECT 0.2190 0.2730 0.3660 0.2870 ;
         RECT 0.3655 0.0920 0.3875 0.1540 ;
         RECT 0.3655 0.1540 0.3875 0.2730 ;
         RECT 0.3655 0.2730 0.3875 0.2870 ;
         RECT 0.2830 0.0510 0.3050 0.0650 ;
         RECT 0.2830 0.0650 0.3050 0.1670 ;
         RECT 0.2935 0.0510 0.3155 0.0650 ;
        RECT 0.3060 0.0510 0.5790 0.0650 ;
        RECT 0.3060 0.3140 0.5790 0.3380 ;
         RECT 0.5770 0.0510 0.5990 0.0650 ;
         RECT 0.5770 0.0650 0.5990 0.1670 ;
         RECT 0.5770 0.1670 0.5990 0.3140 ;
         RECT 0.5770 0.3140 0.5990 0.3380 ;
  END
END CLKGATETST_X1

MACRO DFFRNQ_X1
  CLASS core ;
  FOREIGN DFFRNQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 1.092 BY 0.384 ;

  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 0.149 0.121 0.171 0.263 ;  
    END
  END D

  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
      RECT 0.462 0.156 0.744 0.180 ;  
      RECT 0.744 0.156 0.870 0.180 ;  
    END
  END RN

  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
      RECT 0.021 0.128 0.043 0.256 ;  
    END
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT 1.045 0.032 1.067 0.352 ;  
    END
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT -0.007 0.370 0.093 0.398 ;
      RECT 0.093 0.370 0.135 0.398 ;
      RECT 0.135 0.370 0.219 0.398 ;
      RECT 0.219 0.370 0.261 0.398 ;
      RECT 0.261 0.370 0.345 0.398 ;
      RECT 0.345 0.370 0.534 0.398 ;
      RECT 0.534 0.370 0.597 0.398 ;
      RECT 0.597 0.370 0.639 0.398 ;
      RECT 0.639 0.370 0.723 0.398 ;
      RECT 0.723 0.370 0.780 0.398 ;
      RECT 0.780 0.370 0.977 0.398 ;
      RECT 0.977 0.370 1.099 0.398 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT -0.007 -0.014 1.099 0.014 ;
    END
  END VSS

  OBS
    LAYER MINT1 ;
      RECT 0.0958125 0.137812 0.744125 0.156187 ;
      RECT 0.0538125 0.347813 0.744125 0.366187 ;
    LAYER MINT1 ;
      RECT 0.0958125 0.137812 0.744125 0.156187 ;
      RECT 0.0538125 0.347813 0.744125 0.366187 ;
    LAYER M1 ;
      RECT 0.117 0.036 0.135 0.348 ;
      RECT 0.201 0.036 0.219 0.348 ;
      RECT 0.348 0.312 0.534 0.340 ;
      RECT 0.285 0.051 0.303 0.065 ;
      RECT 0.285 0.065 0.303 0.219 ;
      RECT 0.285 0.219 0.303 0.335 ;
      RECT 0.303 0.051 0.525 0.065 ;
      RECT 0.525 0.051 0.543 0.065 ;
      RECT 0.525 0.065 0.543 0.219 ;
      RECT 0.378 0.165 0.396 0.253 ;
      RECT 0.378 0.253 0.396 0.267 ;
      RECT 0.396 0.253 0.579 0.267 ;
      RECT 0.579 0.036 0.597 0.165 ;
      RECT 0.579 0.165 0.597 0.253 ;
      RECT 0.579 0.253 0.579 0.267 ;
      RECT 0.579 0.267 0.597 0.336 ;
      RECT 0.663 0.051 0.681 0.065 ;
      RECT 0.663 0.065 0.681 0.183 ;
      RECT 0.663 0.183 0.681 0.335 ;
      RECT 0.681 0.051 0.876 0.065 ;
      RECT 0.876 0.051 0.894 0.065 ;
      RECT 0.876 0.065 0.894 0.183 ;
      RECT 0.803 0.197 0.822 0.319 ;
      RECT 0.803 0.319 0.822 0.333 ;
      RECT 0.822 0.319 0.957 0.333 ;
      RECT 0.957 0.036 0.975 0.066 ;
      RECT 0.957 0.066 0.975 0.197 ;
      RECT 0.957 0.197 0.975 0.319 ;
      RECT 0.957 0.319 0.975 0.333 ;
      RECT 0.975 0.066 0.977 0.197 ;
      RECT 0.975 0.197 0.977 0.319 ;
      RECT 0.975 0.319 0.977 0.333 ;
      RECT 0.032 0.042 0.052 0.070 ;
      RECT 0.032 0.070 0.052 0.084 ;
      RECT 0.032 0.283 0.052 0.303 ;
      RECT 0.032 0.303 0.052 0.343 ;
      RECT 0.052 0.070 0.075 0.084 ;
      RECT 0.052 0.283 0.075 0.303 ;
      RECT 0.075 0.070 0.093 0.084 ;
      RECT 0.075 0.084 0.093 0.283 ;
      RECT 0.075 0.283 0.093 0.303 ;
      RECT 0.243 0.097 0.261 0.247 ;
      RECT 0.327 0.201 0.345 0.287 ;
      RECT 0.345 0.097 0.366 0.147 ;
      RECT 0.483 0.129 0.501 0.219 ;
      RECT 0.621 0.137 0.639 0.289 ;
      RECT 0.705 0.087 0.723 0.158 ;
      RECT 0.705 0.230 0.723 0.311 ;
      RECT 0.759 0.083 0.780 0.343 ;
      RECT 0.831 0.087 0.849 0.159 ;
    LAYER V1 ;
      RECT 0.075 0.265 0.093 0.279 ;
      RECT 0.117 0.105 0.135 0.119 ;
      RECT 0.243 0.105 0.261 0.119 ;
      RECT 0.327 0.265 0.345 0.279 ;
      RECT 0.348 0.105 0.366 0.119 ;
      RECT 0.483 0.137 0.501 0.151 ;
      RECT 0.621 0.265 0.639 0.279 ;
      RECT 0.705 0.105 0.723 0.119 ;
      RECT 0.705 0.265 0.723 0.279 ;
      RECT 0.831 0.137 0.849 0.151 ;
    LAYER M1 ;
      RECT 0.117 0.036 0.135 0.348 ;
      RECT 0.201 0.036 0.219 0.348 ;
      RECT 0.348 0.312 0.534 0.340 ;
      RECT 0.285 0.051 0.303 0.065 ;
      RECT 0.285 0.065 0.303 0.219 ;
      RECT 0.285 0.219 0.303 0.335 ;
      RECT 0.303 0.051 0.525 0.065 ;
      RECT 0.525 0.051 0.543 0.065 ;
      RECT 0.525 0.065 0.543 0.219 ;
      RECT 0.378 0.165 0.396 0.253 ;
      RECT 0.378 0.253 0.396 0.267 ;
      RECT 0.396 0.253 0.579 0.267 ;
      RECT 0.579 0.036 0.597 0.165 ;
      RECT 0.579 0.165 0.597 0.253 ;
      RECT 0.579 0.253 0.579 0.267 ;
      RECT 0.579 0.267 0.579 0.336 ;
      RECT 0.663 0.051 0.681 0.065 ;
      RECT 0.663 0.065 0.681 0.183 ;
      RECT 0.663 0.183 0.681 0.335 ;
      RECT 0.681 0.051 0.876 0.065 ;
      RECT 0.876 0.051 0.894 0.065 ;
      RECT 0.876 0.065 0.894 0.183 ;
      RECT 0.803 0.197 0.822 0.319 ;
      RECT 0.803 0.319 0.822 0.333 ;
      RECT 0.822 0.319 0.957 0.333 ;
      RECT 0.957 0.036 0.975 0.066 ;
      RECT 0.957 0.066 0.975 0.197 ;
      RECT 0.957 0.197 0.975 0.319 ;
      RECT 0.957 0.319 0.975 0.333 ;
      RECT 0.975 0.066 0.977 0.197 ;
      RECT 0.975 0.197 0.977 0.319 ;
      RECT 0.975 0.319 0.977 0.333 ;
      RECT 0.032 0.042 0.052 0.070 ;
      RECT 0.032 0.070 0.052 0.084 ;
      RECT 0.032 0.283 0.052 0.303 ;
      RECT 0.032 0.303 0.052 0.343 ;
      RECT 0.052 0.070 0.075 0.084 ;
      RECT 0.052 0.283 0.075 0.303 ;
      RECT 0.075 0.070 0.093 0.084 ;
      RECT 0.075 0.084 0.093 0.283 ;
      RECT 0.075 0.283 0.093 0.303 ;
      RECT 0.243 0.097 0.261 0.247 ;
      RECT 0.327 0.201 0.345 0.287 ;
      RECT 0.345 0.097 0.366 0.147 ;
      RECT 0.483 0.129 0.501 0.219 ;
      RECT 0.621 0.137 0.639 0.289 ;
      RECT 0.705 0.087 0.723 0.158 ;
      RECT 0.705 0.230 0.723 0.311 ;
      RECT 0.759 0.083 0.780 0.343 ;
      RECT 0.831 0.087 0.849 0.159 ;
  END
END DFFRNQ_X1

MACRO DFFSNQ_X1
  CLASS core ;
  FOREIGN DFFSNQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 1.0920 BY 0.3840 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1570 0.1210 0.1790 0.2630 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
         RECT 0.4740 0.1320 0.7440 0.1560 ;
         RECT 0.7440 0.1320 0.8700 0.1560 ;
    END
  END SN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1280 0.0530 0.2560 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 1.0390 0.0320 1.0610 0.3520 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.0930 0.3980 ;
        RECT 0.0930 0.3700 0.1350 0.3980 ;
        RECT 0.1350 0.3700 0.2190 0.3980 ;
        RECT 0.2190 0.3700 0.2610 0.3980 ;
        RECT 0.2610 0.3700 0.3450 0.3980 ;
         RECT 0.3435 0.3700 0.3655 0.3980 ;
        RECT 0.3640 0.3700 0.5970 0.3980 ;
        RECT 0.5970 0.3700 0.6390 0.3980 ;
        RECT 0.6390 0.3700 0.7260 0.3980 ;
        RECT 0.7260 0.3700 0.9120 0.3980 ;
        RECT 0.9120 0.3700 0.9760 0.3980 ;
        RECT 0.9760 0.3700 1.0990 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 1.0990 0.0140 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
         RECT 0.0960 0.1000 0.7440 0.1240 ;
         RECT 0.0540 0.2600 0.7440 0.2840 ;
      LAYER MINT1 ;
         RECT 0.0960 0.1000 0.7440 0.1240 ;
         RECT 0.0540 0.2600 0.7440 0.2840 ;
      LAYER M1 ;
         RECT 0.1150 0.0360 0.1370 0.3480 ;
         RECT 0.1990 0.0360 0.2210 0.3480 ;
         RECT 0.2830 0.0610 0.3050 0.0750 ;
         RECT 0.2830 0.0750 0.3050 0.1830 ;
         RECT 0.2830 0.1830 0.3050 0.3350 ;
        RECT 0.3030 0.0610 0.5370 0.0750 ;
         RECT 0.5350 0.0610 0.5570 0.0750 ;
         RECT 0.5350 0.0750 0.5570 0.1830 ;
         RECT 0.6190 0.1370 0.6410 0.2870 ;
         RECT 0.7045 0.0970 0.7265 0.1620 ;
         RECT 0.7045 0.1960 0.7265 0.2970 ;
         RECT 0.8290 0.0930 0.8510 0.1590 ;
         RECT 0.7870 0.1970 0.8090 0.2870 ;
         RECT 0.7870 0.2870 0.8090 0.3010 ;
        RECT 0.8070 0.2870 0.9570 0.3010 ;
         RECT 0.9550 0.0360 0.9770 0.0660 ;
         RECT 0.9550 0.0660 0.9770 0.1970 ;
         RECT 0.9550 0.1970 0.9770 0.2870 ;
         RECT 0.9550 0.2870 0.9770 0.3010 ;
         RECT 0.9645 0.0660 0.9865 0.1970 ;
         RECT 0.9645 0.1970 0.9865 0.2870 ;
         RECT 0.9645 0.2870 0.9865 0.3010 ;
         RECT 0.0200 0.0410 0.0420 0.0690 ;
         RECT 0.0200 0.0690 0.0420 0.0880 ;
         RECT 0.0310 0.0410 0.0530 0.0690 ;
         RECT 0.0310 0.0690 0.0530 0.0880 ;
         RECT 0.0310 0.2830 0.0530 0.3030 ;
         RECT 0.0310 0.3030 0.0530 0.3430 ;
         RECT 0.0420 0.0410 0.0640 0.0690 ;
         RECT 0.0420 0.0690 0.0640 0.0880 ;
         RECT 0.0420 0.2830 0.0640 0.3030 ;
         RECT 0.0535 0.0690 0.0755 0.0880 ;
         RECT 0.0535 0.2830 0.0755 0.3030 ;
         RECT 0.0730 0.0690 0.0950 0.0880 ;
         RECT 0.0730 0.0880 0.0950 0.2830 ;
         RECT 0.0730 0.2830 0.0950 0.3030 ;
         RECT 0.2410 0.0970 0.2630 0.2470 ;
         RECT 0.3250 0.2010 0.3470 0.2950 ;
         RECT 0.3435 0.0970 0.3655 0.1520 ;
         RECT 0.4930 0.1290 0.5150 0.1830 ;
         RECT 0.3970 0.1370 0.4190 0.2870 ;
         RECT 0.3970 0.2870 0.4190 0.3010 ;
        RECT 0.4170 0.2870 0.5760 0.3010 ;
         RECT 0.5665 0.2870 0.5885 0.3010 ;
         RECT 0.5665 0.3010 0.5885 0.3430 ;
         RECT 0.5770 0.0480 0.5990 0.1370 ;
         RECT 0.5770 0.1370 0.5990 0.2870 ;
         RECT 0.5770 0.2870 0.5990 0.3010 ;
         RECT 0.5770 0.3010 0.5990 0.3430 ;
         RECT 0.6610 0.0570 0.6830 0.0710 ;
         RECT 0.6610 0.0710 0.6830 0.1830 ;
         RECT 0.6610 0.1830 0.6830 0.3360 ;
        RECT 0.6810 0.0570 0.8870 0.0710 ;
         RECT 0.8855 0.0570 0.9075 0.0710 ;
         RECT 0.8855 0.0710 0.9075 0.1830 ;
        RECT 0.7260 0.3190 0.9120 0.3330 ;
      LAYER V1 ;
        RECT 0.0750 0.2650 0.0930 0.2790 ;
        RECT 0.1170 0.1050 0.1350 0.1190 ;
        RECT 0.2430 0.1050 0.2610 0.1190 ;
        RECT 0.3270 0.2650 0.3450 0.2790 ;
        RECT 0.3450 0.1050 0.3640 0.1190 ;
        RECT 0.4950 0.1370 0.5130 0.1510 ;
        RECT 0.6210 0.2650 0.6390 0.2790 ;
        RECT 0.7050 0.1050 0.7230 0.1190 ;
        RECT 0.7050 0.2650 0.7230 0.2790 ;
        RECT 0.8310 0.1370 0.8490 0.1510 ;
      LAYER M1 ;
         RECT 0.1150 0.0360 0.1370 0.3480 ;
         RECT 0.1990 0.0360 0.2210 0.3480 ;
         RECT 0.2830 0.0610 0.3050 0.0750 ;
         RECT 0.2830 0.0750 0.3050 0.1830 ;
         RECT 0.2830 0.1830 0.3050 0.3350 ;
        RECT 0.3030 0.0610 0.5370 0.0750 ;
         RECT 0.5350 0.0610 0.5570 0.0750 ;
         RECT 0.5350 0.0750 0.5570 0.1830 ;
         RECT 0.6190 0.1370 0.6410 0.2870 ;
         RECT 0.7045 0.0970 0.7265 0.1620 ;
         RECT 0.7045 0.1960 0.7265 0.2970 ;
         RECT 0.8290 0.0930 0.8510 0.1590 ;
         RECT 0.7870 0.1970 0.8090 0.2870 ;
         RECT 0.7870 0.2870 0.8090 0.3010 ;
        RECT 0.8070 0.2870 0.9570 0.3010 ;
         RECT 0.9550 0.0360 0.9770 0.0660 ;
         RECT 0.9550 0.0660 0.9770 0.1970 ;
         RECT 0.9550 0.1970 0.9770 0.2870 ;
         RECT 0.9550 0.2870 0.9770 0.3010 ;
         RECT 0.9645 0.0660 0.9865 0.1970 ;
         RECT 0.9645 0.1970 0.9865 0.2870 ;
         RECT 0.9645 0.2870 0.9865 0.3010 ;
         RECT 0.0200 0.0410 0.0420 0.0690 ;
         RECT 0.0200 0.0690 0.0420 0.0880 ;
         RECT 0.0310 0.0410 0.0530 0.0690 ;
         RECT 0.0310 0.0690 0.0530 0.0880 ;
         RECT 0.0310 0.2830 0.0530 0.3030 ;
         RECT 0.0310 0.3030 0.0530 0.3430 ;
         RECT 0.0420 0.0410 0.0640 0.0690 ;
         RECT 0.0420 0.0690 0.0640 0.0880 ;
         RECT 0.0420 0.2830 0.0640 0.3030 ;
         RECT 0.0535 0.0690 0.0755 0.0880 ;
         RECT 0.0535 0.2830 0.0755 0.3030 ;
         RECT 0.0730 0.0690 0.0950 0.0880 ;
         RECT 0.0730 0.0880 0.0950 0.2830 ;
         RECT 0.0730 0.2830 0.0950 0.3030 ;
         RECT 0.2410 0.0970 0.2630 0.2470 ;
         RECT 0.3250 0.2010 0.3470 0.2950 ;
         RECT 0.3435 0.0970 0.3655 0.1520 ;
         RECT 0.4930 0.1290 0.5150 0.1830 ;
         RECT 0.3970 0.1370 0.4190 0.2870 ;
         RECT 0.3970 0.2870 0.4190 0.3010 ;
        RECT 0.4170 0.2870 0.5760 0.3010 ;
         RECT 0.5665 0.2870 0.5885 0.3010 ;
         RECT 0.5665 0.3010 0.5885 0.3430 ;
         RECT 0.5770 0.0480 0.5990 0.1370 ;
         RECT 0.5770 0.1370 0.5990 0.2870 ;
         RECT 0.5770 0.2870 0.5990 0.3010 ;
         RECT 0.5770 0.3010 0.5990 0.3430 ;
         RECT 0.6610 0.0570 0.6830 0.0710 ;
         RECT 0.6610 0.0710 0.6830 0.1830 ;
         RECT 0.6610 0.1830 0.6830 0.3360 ;
        RECT 0.6810 0.0570 0.8870 0.0710 ;
         RECT 0.8855 0.0570 0.9075 0.0710 ;
         RECT 0.8855 0.0710 0.9075 0.1830 ;
        RECT 0.7260 0.3190 0.9120 0.3330 ;
  END
END DFFSNQ_X1

MACRO FA_X1
  CLASS core ;
  FOREIGN FA_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 1.0080 BY 0.3840 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
         RECT 0.1380 0.2280 0.7210 0.2520 ;
      LAYER V1 ;
        RECT 0.4300 0.2330 0.4490 0.2470 ;
        RECT 0.6810 0.2330 0.7000 0.2470 ;
      LAYER M1 ;
         RECT 0.4285 0.2010 0.4505 0.2630 ;
        RECT 0.6810 0.1370 0.7050 0.2630 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
         RECT 0.1800 0.1320 0.5180 0.1560 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
         RECT 0.0960 0.1000 0.8280 0.1240 ;
      LAYER V1 ;
        RECT 0.1170 0.1050 0.1350 0.1190 ;
        RECT 0.3810 0.1050 0.3990 0.1190 ;
        RECT 0.7890 0.1050 0.8070 0.1190 ;
      LAYER M1 ;
         RECT 0.1150 0.0970 0.1370 0.2950 ;
         RECT 0.3790 0.0970 0.4010 0.1830 ;
         RECT 0.7870 0.0890 0.8090 0.1830 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.9550 0.0570 0.9770 0.3270 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.5350 0.1030 0.5570 0.3200 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.0930 0.3980 ;
        RECT 0.0930 0.3700 0.1770 0.3980 ;
        RECT 0.1770 0.3700 0.2190 0.3980 ;
        RECT 0.2190 0.3700 0.4300 0.3980 ;
        RECT 0.4300 0.3700 0.5030 0.3980 ;
        RECT 0.5030 0.3700 0.6810 0.3980 ;
        RECT 0.6810 0.3700 0.7110 0.3980 ;
        RECT 0.7110 0.3700 0.7650 0.3980 ;
        RECT 0.7650 0.3700 0.8460 0.3980 ;
        RECT 0.8460 0.3700 0.8910 0.3980 ;
        RECT 0.8910 0.3700 1.0150 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 1.0150 0.0140 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
         RECT 0.0540 0.1960 0.8670 0.2200 ;
         RECT 0.2640 0.1640 0.9120 0.1880 ;
      LAYER MINT1 ;
         RECT 0.0540 0.1960 0.8670 0.2200 ;
         RECT 0.2640 0.1640 0.9120 0.1880 ;
      LAYER M1 ;
        RECT 0.0180 0.0890 0.0430 0.1690 ;
        RECT 0.0180 0.1690 0.0430 0.1830 ;
        RECT 0.0430 0.1690 0.0680 0.1830 ;
        RECT 0.0680 0.1690 0.0930 0.1830 ;
        RECT 0.0680 0.1830 0.0930 0.2310 ;
         RECT 0.1570 0.1370 0.1790 0.2950 ;
        RECT 0.2780 0.1370 0.3030 0.2540 ;
        RECT 0.2430 0.0480 0.4060 0.0680 ;
         RECT 0.2425 0.2880 0.2645 0.3020 ;
         RECT 0.2425 0.3020 0.2645 0.3490 ;
        RECT 0.2640 0.2880 0.4090 0.3020 ;
         RECT 0.4085 0.2880 0.4305 0.3020 ;
         RECT 0.4085 0.3020 0.4305 0.3490 ;
         RECT 0.4085 0.3490 0.4305 0.3520 ;
        RECT 0.4780 0.1220 0.5030 0.2320 ;
         RECT 0.5770 0.0970 0.5990 0.1830 ;
         RECT 0.5770 0.2810 0.5990 0.2950 ;
         RECT 0.5770 0.2950 0.5990 0.3480 ;
        RECT 0.5970 0.2810 0.6630 0.2950 ;
         RECT 0.6610 0.2810 0.6830 0.2950 ;
         RECT 0.6610 0.2950 0.6830 0.3480 ;
         RECT 0.7450 0.0360 0.7670 0.3480 ;
         RECT 0.8255 0.1930 0.8475 0.2950 ;
         RECT 0.1990 0.0480 0.2210 0.3360 ;
         RECT 0.3250 0.1370 0.3470 0.2540 ;
        RECT 0.6210 0.1370 0.6460 0.2470 ;
        RECT 0.5550 0.0500 0.7110 0.0660 ;
         RECT 0.8710 0.1370 0.8930 0.2630 ;
      LAYER V1 ;
        RECT 0.0750 0.2010 0.0930 0.2150 ;
        RECT 0.1590 0.2330 0.1770 0.2470 ;
        RECT 0.2010 0.1370 0.2190 0.1510 ;
        RECT 0.2850 0.1690 0.3030 0.1830 ;
        RECT 0.3270 0.2010 0.3450 0.2150 ;
        RECT 0.4780 0.1370 0.4970 0.1510 ;
        RECT 0.5790 0.1050 0.5970 0.1190 ;
        RECT 0.6270 0.2010 0.6460 0.2150 ;
        RECT 0.7470 0.1690 0.7650 0.1830 ;
        RECT 0.8270 0.2010 0.8460 0.2150 ;
        RECT 0.8730 0.1690 0.8910 0.1830 ;
      LAYER M1 ;
        RECT 0.0180 0.0890 0.0430 0.1690 ;
        RECT 0.0180 0.1690 0.0430 0.1830 ;
        RECT 0.0430 0.1690 0.0680 0.1830 ;
        RECT 0.0680 0.1690 0.0930 0.1830 ;
        RECT 0.0680 0.1830 0.0930 0.2310 ;
         RECT 0.1570 0.1370 0.1790 0.2950 ;
        RECT 0.2780 0.1370 0.3030 0.2540 ;
        RECT 0.2430 0.0480 0.4060 0.0680 ;
         RECT 0.2425 0.2880 0.2645 0.3020 ;
         RECT 0.2425 0.3020 0.2645 0.3490 ;
        RECT 0.2640 0.2880 0.4090 0.3020 ;
         RECT 0.4085 0.2880 0.4305 0.3020 ;
         RECT 0.4085 0.3020 0.4305 0.3490 ;
         RECT 0.4085 0.3490 0.4305 0.3520 ;
        RECT 0.4780 0.1220 0.5030 0.2320 ;
         RECT 0.5770 0.0970 0.5990 0.1830 ;
         RECT 0.5770 0.2810 0.5990 0.2950 ;
         RECT 0.5770 0.2950 0.5990 0.3480 ;
        RECT 0.5970 0.2810 0.6630 0.2950 ;
         RECT 0.6610 0.2810 0.6830 0.2950 ;
         RECT 0.6610 0.2950 0.6830 0.3480 ;
         RECT 0.7450 0.0360 0.7670 0.3480 ;
         RECT 0.8255 0.1930 0.8475 0.2950 ;
         RECT 0.1990 0.0480 0.2210 0.3360 ;
         RECT 0.3250 0.1370 0.3470 0.2540 ;
        RECT 0.6210 0.1370 0.6460 0.2470 ;
        RECT 0.5550 0.0500 0.7110 0.0660 ;
         RECT 0.8710 0.1370 0.8930 0.2630 ;
  END
END FA_X1

MACRO FILLTIE
  CLASS core ;
  FOREIGN FILLTIE 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.3780 BY 0.3840 ;
  OBS
      LAYER M1 ;
        RECT 0.0010 0.0010 0.3860 0.0140 ;
        RECT 0.0010 0.3700 0.3860 0.3980 ;
      LAYER M1 ;
        RECT 0.0010 0.0010 0.3860 0.0140 ;
        RECT 0.0010 0.3700 0.3860 0.3980 ;
  END
END FILLTIE

MACRO FILL_X1
  CLASS core ;
  FOREIGN FILL_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.0840 BY 0.3840 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.0910 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.0910 0.0140 ;
    END
  END VSS
END FILL_X1

MACRO FILL_X2
  CLASS core ;
  FOREIGN FILL_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.1260 BY 0.3840 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.1330 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.1330 0.0140 ;
    END
  END VSS
END FILL_X2

MACRO FILL_X4
  CLASS core ;
  FOREIGN FILL_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.2100 BY 0.3840 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.2170 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.2170 0.0140 ;
    END
  END VSS
END FILL_X4

MACRO FILL_X8
  CLASS core ;
  FOREIGN FILL_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.3780 BY 0.3840 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.3850 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.3850 0.0140 ;
    END
  END VSS
END FILL_X8

MACRO FILL_X16
  CLASS core ;
  FOREIGN FILL_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.7140 BY 0.3840 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.7210 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.7210 0.0140 ;
    END
  END VSS
END FILL_X16

MACRO HA_X1
  CLASS core ;
  FOREIGN HA_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.5460 BY 0.3840 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1570 0.1370 0.1790 0.2780 ;
         RECT 0.1570 0.2780 0.1790 0.2920 ;
        RECT 0.1770 0.2780 0.2850 0.2920 ;
         RECT 0.2830 0.1370 0.3050 0.2780 ;
         RECT 0.2830 0.2780 0.3050 0.2920 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1990 0.1280 0.2210 0.2560 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.0410 0.0530 0.3190 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.4930 0.0900 0.5150 0.3190 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.3910 0.3980 ;
        RECT 0.3910 0.3700 0.4330 0.3980 ;
        RECT 0.4330 0.3700 0.5530 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.5530 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.2220 0.0510 0.4080 0.0650 ;
        RECT 0.2660 0.0920 0.3270 0.1080 ;
         RECT 0.3265 0.0920 0.3485 0.1080 ;
         RECT 0.3265 0.1080 0.3485 0.2310 ;
         RECT 0.3265 0.2310 0.3485 0.3010 ;
        RECT 0.3480 0.0920 0.4150 0.1080 ;
         RECT 0.4130 0.0920 0.4350 0.1080 ;
         RECT 0.4130 0.1080 0.4350 0.2310 ;
         RECT 0.0730 0.0830 0.0950 0.0990 ;
         RECT 0.0730 0.0990 0.0950 0.1370 ;
         RECT 0.0730 0.1370 0.0950 0.3190 ;
         RECT 0.0730 0.3190 0.0950 0.3330 ;
        RECT 0.0930 0.0830 0.2430 0.0990 ;
        RECT 0.0930 0.3190 0.2430 0.3330 ;
        RECT 0.2430 0.3190 0.3710 0.3330 ;
         RECT 0.3700 0.1370 0.3920 0.3190 ;
         RECT 0.3700 0.3190 0.3920 0.3330 ;
      LAYER M1 ;
        RECT 0.2220 0.0510 0.4080 0.0650 ;
        RECT 0.2660 0.0920 0.3270 0.1080 ;
         RECT 0.3265 0.0920 0.3485 0.1080 ;
         RECT 0.3265 0.1080 0.3485 0.2310 ;
         RECT 0.3265 0.2310 0.3485 0.3010 ;
        RECT 0.3480 0.0920 0.4150 0.1080 ;
         RECT 0.4130 0.0920 0.4350 0.1080 ;
         RECT 0.4130 0.1080 0.4350 0.2310 ;
         RECT 0.0730 0.0830 0.0950 0.0990 ;
         RECT 0.0730 0.0990 0.0950 0.1370 ;
         RECT 0.0730 0.1370 0.0950 0.3190 ;
         RECT 0.0730 0.3190 0.0950 0.3330 ;
        RECT 0.0930 0.0830 0.2430 0.0990 ;
        RECT 0.0930 0.3190 0.2430 0.3330 ;
        RECT 0.2430 0.3190 0.3710 0.3330 ;
         RECT 0.3700 0.1370 0.3920 0.3190 ;
         RECT 0.3700 0.3190 0.3920 0.3330 ;
  END
END HA_X1

MACRO INV_X1
  CLASS core ;
  FOREIGN INV_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.1260 BY 0.3840 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.0960 0.0530 0.2880 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.0570 0.0950 0.3200 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.1330 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.1330 0.0140 ;
    END
  END VSS
END INV_X1

MACRO INV_X2
  CLASS core ;
  FOREIGN INV_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.1680 BY 0.3840 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.0960 0.0530 0.2880 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.0650 0.0950 0.2880 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.1750 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.1750 0.0140 ;
    END
  END VSS
END INV_X2

MACRO INV_X4
  CLASS core ;
  FOREIGN INV_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.2520 BY 0.3840 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1280 0.0530 0.1840 ;
         RECT 0.0310 0.1840 0.0530 0.1980 ;
         RECT 0.0310 0.1980 0.0530 0.2560 ;
        RECT 0.0520 0.1840 0.1560 0.1980 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0220 0.0710 0.0440 0.1000 ;
        RECT 0.0390 0.0710 0.2010 0.1000 ;
        RECT 0.0390 0.2840 0.2010 0.3130 ;
         RECT 0.1990 0.0710 0.2210 0.1000 ;
         RECT 0.1990 0.1000 0.2210 0.2840 ;
         RECT 0.1990 0.2840 0.2210 0.3130 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.2590 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.2590 0.0140 ;
    END
  END VSS
END INV_X4

MACRO INV_X8
  CLASS core ;
  FOREIGN INV_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.4200 BY 0.3840 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.0970 0.0950 0.1980 ;
         RECT 0.0730 0.1980 0.0950 0.2280 ;
         RECT 0.0730 0.2280 0.0950 0.2880 ;
        RECT 0.0930 0.1980 0.3030 0.2280 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0200 0.3160 0.0420 0.3300 ;
        RECT 0.0350 0.0550 0.3660 0.0690 ;
        RECT 0.0350 0.3160 0.3660 0.3300 ;
        RECT 0.3660 0.0550 0.3900 0.0690 ;
        RECT 0.3660 0.0690 0.3900 0.3160 ;
        RECT 0.3660 0.3160 0.3900 0.3300 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.4270 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.4270 0.0140 ;
    END
  END VSS
END INV_X8

MACRO INV_X12
  CLASS core ;
  FOREIGN INV_X12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.5880 BY 0.3840 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.0960 0.0950 0.1840 ;
         RECT 0.0730 0.1840 0.0950 0.1980 ;
         RECT 0.0730 0.1980 0.0950 0.2880 ;
        RECT 0.0930 0.1840 0.4500 0.1980 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.0350 0.0510 0.5330 0.0650 ;
        RECT 0.0350 0.3180 0.5330 0.3340 ;
        RECT 0.5330 0.0510 0.5580 0.0650 ;
        RECT 0.5330 0.0650 0.5580 0.3180 ;
        RECT 0.5330 0.3180 0.5580 0.3340 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.5950 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.5950 0.0140 ;
    END
  END VSS
END INV_X12

MACRO INV_X16
  CLASS core ;
  FOREIGN INV_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.7560 BY 0.3840 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1280 0.0530 0.1850 ;
         RECT 0.0310 0.1850 0.0530 0.1990 ;
         RECT 0.0310 0.1990 0.0530 0.2810 ;
        RECT 0.0510 0.1850 0.6180 0.1990 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.7020 0.3980 ;
        RECT 0.7020 0.3700 0.7630 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.7630 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.0350 0.0500 0.6810 0.0660 ;
        RECT 0.0350 0.3110 0.6810 0.3400 ;
         RECT 0.6805 0.0500 0.7025 0.0660 ;
         RECT 0.6805 0.0660 0.7025 0.3110 ;
         RECT 0.6805 0.3110 0.7025 0.3400 ;
      LAYER M1 ;
        RECT 0.0350 0.0500 0.6810 0.0660 ;
        RECT 0.0350 0.3110 0.6810 0.3400 ;
         RECT 0.6805 0.0500 0.7025 0.0660 ;
         RECT 0.6805 0.0660 0.7025 0.3110 ;
         RECT 0.6805 0.3110 0.7025 0.3400 ;
  END
END INV_X16

MACRO LHQ_X1
  CLASS core ;
  FOREIGN LHQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.5880 BY 0.3840 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1570 0.0800 0.1790 0.2560 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1280 0.0530 0.2560 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.5350 0.0650 0.5570 0.3190 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.5130 0.3980 ;
        RECT 0.5130 0.3700 0.5950 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.5950 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0215 0.2780 0.0435 0.2920 ;
         RECT 0.0215 0.2920 0.0435 0.3520 ;
         RECT 0.0310 0.0320 0.0530 0.0460 ;
         RECT 0.0310 0.0460 0.0530 0.0920 ;
         RECT 0.0310 0.0920 0.0530 0.1060 ;
         RECT 0.0310 0.2780 0.0530 0.2920 ;
         RECT 0.0310 0.2920 0.0530 0.3520 ;
         RECT 0.0405 0.0320 0.0625 0.0460 ;
         RECT 0.0405 0.0920 0.0625 0.1060 ;
         RECT 0.0405 0.2780 0.0625 0.2920 ;
         RECT 0.0405 0.2920 0.0625 0.3520 ;
        RECT 0.0520 0.0320 0.0750 0.0460 ;
        RECT 0.0520 0.0920 0.0750 0.1060 ;
        RECT 0.0520 0.2780 0.0750 0.2920 ;
         RECT 0.0730 0.0320 0.0950 0.0460 ;
         RECT 0.0730 0.0920 0.0950 0.1060 ;
         RECT 0.0730 0.1060 0.0950 0.1610 ;
         RECT 0.0730 0.1610 0.0950 0.1750 ;
         RECT 0.0730 0.1750 0.0950 0.2070 ;
         RECT 0.0730 0.2070 0.0950 0.2780 ;
         RECT 0.0730 0.2780 0.0950 0.2920 ;
        RECT 0.0930 0.0320 0.2130 0.0460 ;
         RECT 0.2110 0.0320 0.2330 0.0460 ;
         RECT 0.2110 0.0460 0.2330 0.0920 ;
         RECT 0.2110 0.0920 0.2330 0.1060 ;
         RECT 0.2110 0.1060 0.2330 0.1610 ;
         RECT 0.2110 0.1610 0.2330 0.1750 ;
         RECT 0.2260 0.1610 0.2480 0.1750 ;
         RECT 0.2410 0.1610 0.2630 0.1750 ;
         RECT 0.2410 0.1750 0.2630 0.2070 ;
         RECT 0.3460 0.0570 0.3680 0.0710 ;
         RECT 0.3460 0.0710 0.3680 0.2470 ;
        RECT 0.3660 0.0570 0.4530 0.0710 ;
         RECT 0.4510 0.0570 0.4730 0.0710 ;
         RECT 0.4510 0.0710 0.4730 0.2470 ;
         RECT 0.4510 0.2470 0.4730 0.2960 ;
         RECT 0.1150 0.0680 0.1370 0.2300 ;
         RECT 0.1150 0.2300 0.1370 0.2780 ;
         RECT 0.1150 0.2780 0.1370 0.2920 ;
        RECT 0.1350 0.2780 0.2010 0.2920 ;
         RECT 0.2010 0.2300 0.2230 0.2780 ;
         RECT 0.2010 0.2780 0.2230 0.2920 ;
        RECT 0.1800 0.3190 0.2550 0.3330 ;
        RECT 0.2550 0.0570 0.3060 0.0860 ;
        RECT 0.2550 0.3190 0.3060 0.3330 ;
         RECT 0.3040 0.0570 0.3260 0.0860 ;
         RECT 0.3040 0.0860 0.3260 0.1530 ;
         RECT 0.3040 0.1530 0.3260 0.3180 ;
         RECT 0.3040 0.3180 0.3260 0.3190 ;
         RECT 0.3040 0.3190 0.3260 0.3330 ;
        RECT 0.3240 0.3180 0.4950 0.3190 ;
        RECT 0.3240 0.3190 0.4950 0.3330 ;
         RECT 0.4930 0.1530 0.5150 0.3180 ;
         RECT 0.4930 0.3180 0.5150 0.3190 ;
         RECT 0.4930 0.3190 0.5150 0.3330 ;
      LAYER M1 ;
         RECT 0.0215 0.2780 0.0435 0.2920 ;
         RECT 0.0215 0.2920 0.0435 0.3520 ;
         RECT 0.0310 0.0320 0.0530 0.0460 ;
         RECT 0.0310 0.0460 0.0530 0.0920 ;
         RECT 0.0310 0.0920 0.0530 0.1060 ;
         RECT 0.0310 0.2780 0.0530 0.2920 ;
         RECT 0.0310 0.2920 0.0530 0.3520 ;
         RECT 0.0405 0.0320 0.0625 0.0460 ;
         RECT 0.0405 0.0920 0.0625 0.1060 ;
         RECT 0.0405 0.2780 0.0625 0.2920 ;
         RECT 0.0405 0.2920 0.0625 0.3520 ;
        RECT 0.0520 0.0320 0.0750 0.0460 ;
        RECT 0.0520 0.0920 0.0750 0.1060 ;
        RECT 0.0520 0.2780 0.0750 0.2920 ;
         RECT 0.0730 0.0320 0.0950 0.0460 ;
         RECT 0.0730 0.0920 0.0950 0.1060 ;
         RECT 0.0730 0.1060 0.0950 0.1610 ;
         RECT 0.0730 0.1610 0.0950 0.1750 ;
         RECT 0.0730 0.1750 0.0950 0.2070 ;
         RECT 0.0730 0.2070 0.0950 0.2780 ;
         RECT 0.0730 0.2780 0.0950 0.2920 ;
        RECT 0.0930 0.0320 0.2130 0.0460 ;
         RECT 0.2110 0.0320 0.2330 0.0460 ;
         RECT 0.2110 0.0460 0.2330 0.0920 ;
         RECT 0.2110 0.0920 0.2330 0.1060 ;
         RECT 0.2110 0.1060 0.2330 0.1610 ;
         RECT 0.2110 0.1610 0.2330 0.1750 ;
         RECT 0.2260 0.1610 0.2480 0.1750 ;
         RECT 0.2410 0.1610 0.2630 0.1750 ;
         RECT 0.2410 0.1750 0.2630 0.2070 ;
         RECT 0.3460 0.0570 0.3680 0.0710 ;
         RECT 0.3460 0.0710 0.3680 0.2470 ;
        RECT 0.3660 0.0570 0.4530 0.0710 ;
         RECT 0.4510 0.0570 0.4730 0.0710 ;
         RECT 0.4510 0.0710 0.4730 0.2470 ;
         RECT 0.4510 0.2470 0.4730 0.2960 ;
         RECT 0.1150 0.0680 0.1370 0.2300 ;
         RECT 0.1150 0.2300 0.1370 0.2780 ;
         RECT 0.1150 0.2780 0.1370 0.2920 ;
        RECT 0.1350 0.2780 0.2010 0.2920 ;
         RECT 0.2010 0.2300 0.2230 0.2780 ;
         RECT 0.2010 0.2780 0.2230 0.2920 ;
        RECT 0.1800 0.3190 0.2550 0.3330 ;
        RECT 0.2550 0.0570 0.3060 0.0860 ;
        RECT 0.2550 0.3190 0.3060 0.3330 ;
         RECT 0.3040 0.0570 0.3260 0.0860 ;
         RECT 0.3040 0.0860 0.3260 0.1530 ;
         RECT 0.3040 0.1530 0.3260 0.3180 ;
         RECT 0.3040 0.3180 0.3260 0.3190 ;
         RECT 0.3040 0.3190 0.3260 0.3330 ;
        RECT 0.3240 0.3180 0.4950 0.3190 ;
        RECT 0.3240 0.3190 0.4950 0.3330 ;
         RECT 0.4930 0.1530 0.5150 0.3180 ;
         RECT 0.4930 0.3180 0.5150 0.3190 ;
         RECT 0.4930 0.3190 0.5150 0.3330 ;
  END
END LHQ_X1

MACRO MUX2_X1
  CLASS core ;
  FOREIGN MUX2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.5460 BY 0.3840 ;
  PIN I0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.3670 0.1210 0.3890 0.2630 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.1280 0.0950 0.2240 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
         RECT 0.0770 0.3240 0.2590 0.3480 ;
      LAYER V1 ;
        RECT 0.0980 0.3290 0.1350 0.3430 ;
      LAYER M1 ;
         RECT 0.0160 0.1210 0.0380 0.3290 ;
         RECT 0.0160 0.3290 0.0380 0.3430 ;
        RECT 0.0360 0.3290 0.1460 0.3430 ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.4510 0.0960 0.4730 0.3190 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.3030 0.3980 ;
        RECT 0.3030 0.3700 0.3450 0.3980 ;
        RECT 0.3450 0.3700 0.5130 0.3980 ;
        RECT 0.5130 0.3700 0.5530 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.5530 0.0140 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
         RECT 0.1800 0.1640 0.3660 0.1880 ;
      LAYER MINT1 ;
         RECT 0.1800 0.1640 0.3660 0.1880 ;
      LAYER M1 ;
         RECT 0.0475 0.0810 0.0695 0.0950 ;
        RECT 0.0650 0.0810 0.1030 0.0950 ;
        RECT 0.0650 0.2460 0.1030 0.2600 ;
        RECT 0.0650 0.2600 0.1030 0.2880 ;
        RECT 0.1030 0.0810 0.2010 0.0950 ;
        RECT 0.1030 0.2460 0.2010 0.2600 ;
         RECT 0.1990 0.0810 0.2210 0.0950 ;
         RECT 0.1990 0.0950 0.2210 0.2460 ;
         RECT 0.1990 0.2460 0.2210 0.2600 ;
        RECT 0.1900 0.3290 0.2850 0.3520 ;
         RECT 0.2830 0.1530 0.3050 0.3290 ;
         RECT 0.2830 0.3290 0.3050 0.3520 ;
         RECT 0.3250 0.1370 0.3470 0.2140 ;
         RECT 0.2410 0.0430 0.2630 0.0730 ;
         RECT 0.2410 0.0730 0.2630 0.2470 ;
         RECT 0.2410 0.2470 0.2630 0.3070 ;
        RECT 0.2610 0.0430 0.4950 0.0730 ;
         RECT 0.4930 0.0430 0.5150 0.0730 ;
         RECT 0.4930 0.0730 0.5150 0.2470 ;
      LAYER V1 ;
        RECT 0.2010 0.1690 0.2190 0.1830 ;
        RECT 0.2010 0.3290 0.2380 0.3430 ;
        RECT 0.3270 0.1690 0.3450 0.1830 ;
      LAYER M1 ;
         RECT 0.0475 0.0810 0.0695 0.0950 ;
        RECT 0.0650 0.0810 0.1030 0.0950 ;
        RECT 0.0650 0.2460 0.1030 0.2600 ;
        RECT 0.0650 0.2600 0.1030 0.2880 ;
        RECT 0.1030 0.0810 0.2010 0.0950 ;
        RECT 0.1030 0.2460 0.2010 0.2600 ;
         RECT 0.1990 0.0810 0.2210 0.0950 ;
         RECT 0.1990 0.0950 0.2210 0.2460 ;
         RECT 0.1990 0.2460 0.2210 0.2600 ;
        RECT 0.1900 0.3290 0.2850 0.3520 ;
         RECT 0.2830 0.1530 0.3050 0.3290 ;
         RECT 0.2830 0.3290 0.3050 0.3520 ;
         RECT 0.3250 0.1370 0.3470 0.2140 ;
         RECT 0.2410 0.0430 0.2630 0.0730 ;
         RECT 0.2410 0.0730 0.2630 0.2470 ;
         RECT 0.2410 0.2470 0.2630 0.3070 ;
        RECT 0.2610 0.0430 0.4950 0.0730 ;
         RECT 0.4930 0.0430 0.5150 0.0730 ;
         RECT 0.4930 0.0730 0.5150 0.2470 ;
  END
END MUX2_X1

MACRO NAND2_X1
  CLASS core ;
  FOREIGN NAND2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.1680 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1150 0.1280 0.1370 0.2870 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1280 0.0530 0.2870 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.0660 0.0950 0.0960 ;
         RECT 0.0730 0.0960 0.0950 0.3190 ;
        RECT 0.0930 0.0660 0.1150 0.0960 ;
         RECT 0.1145 0.0320 0.1365 0.0660 ;
         RECT 0.1145 0.0660 0.1365 0.0960 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.1750 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.1750 0.0140 ;
    END
  END VSS
END NAND2_X1

MACRO NAND2_X2
  CLASS core ;
  FOREIGN NAND2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.2520 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1150 0.1120 0.1370 0.2760 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1370 0.0530 0.3380 ;
         RECT 0.0310 0.3380 0.0530 0.3520 ;
        RECT 0.0510 0.3380 0.2010 0.3520 ;
         RECT 0.1990 0.1370 0.2210 0.3380 ;
         RECT 0.1990 0.3380 0.2210 0.3520 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.0620 0.0950 0.0900 ;
         RECT 0.0730 0.0900 0.0950 0.2120 ;
         RECT 0.0730 0.2120 0.0950 0.2980 ;
         RECT 0.0730 0.2980 0.0950 0.3200 ;
        RECT 0.0930 0.0620 0.1590 0.0900 ;
        RECT 0.0930 0.2980 0.1590 0.3200 ;
         RECT 0.1570 0.0620 0.1790 0.0900 ;
         RECT 0.1570 0.2120 0.1790 0.2980 ;
         RECT 0.1570 0.2980 0.1790 0.3200 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.2590 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.2590 0.0140 ;
    END
  END VSS
END NAND2_X2

MACRO NAND3_X1
  CLASS core ;
  FOREIGN NAND3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.2520 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1570 0.1600 0.1790 0.2240 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1150 0.1280 0.1370 0.2560 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1080 0.0530 0.2870 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.0410 0.0950 0.0550 ;
         RECT 0.0730 0.0550 0.0950 0.1280 ;
         RECT 0.0730 0.1280 0.0950 0.2560 ;
         RECT 0.0730 0.2560 0.0950 0.3380 ;
         RECT 0.0730 0.3380 0.0950 0.3520 ;
        RECT 0.0930 0.0410 0.1590 0.0550 ;
        RECT 0.0930 0.3380 0.1590 0.3520 ;
        RECT 0.1590 0.0320 0.1990 0.0410 ;
        RECT 0.1590 0.0410 0.1990 0.0550 ;
        RECT 0.1590 0.3380 0.1990 0.3520 ;
         RECT 0.1890 0.0320 0.2110 0.0410 ;
         RECT 0.1890 0.0410 0.2110 0.0550 ;
         RECT 0.1890 0.0550 0.2110 0.1280 ;
         RECT 0.1890 0.3380 0.2110 0.3520 ;
         RECT 0.1990 0.0320 0.2210 0.0410 ;
         RECT 0.1990 0.0410 0.2210 0.0550 ;
         RECT 0.1990 0.0550 0.2210 0.1280 ;
         RECT 0.1990 0.2560 0.2210 0.3380 ;
         RECT 0.1990 0.3380 0.2210 0.3520 ;
         RECT 0.2085 0.0320 0.2305 0.0410 ;
         RECT 0.2085 0.0410 0.2305 0.0550 ;
         RECT 0.2085 0.0550 0.2305 0.1280 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.2590 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.2590 0.0140 ;
    END
  END VSS
END NAND3_X1

MACRO NAND3_X2
  CLASS core ;
  FOREIGN NAND3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.3780 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.3250 0.1600 0.3470 0.2560 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1980 0.1240 0.2220 0.2560 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.1280 0.0950 0.2560 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.0180 0.2840 0.2400 0.3130 ;
        RECT 0.2400 0.2840 0.2850 0.3130 ;
         RECT 0.2830 0.0930 0.3050 0.2840 ;
         RECT 0.2830 0.2840 0.3050 0.3130 ;
         RECT 0.3025 0.2840 0.3245 0.3130 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.2400 0.3980 ;
        RECT 0.2400 0.3700 0.3450 0.3980 ;
        RECT 0.3450 0.3700 0.3850 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.3850 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.1380 0.0560 0.3270 0.0700 ;
         RECT 0.3250 0.0560 0.3470 0.0700 ;
         RECT 0.3250 0.0700 0.3470 0.1120 ;
        RECT 0.0330 0.0880 0.2400 0.1040 ;
      LAYER M1 ;
        RECT 0.1380 0.0560 0.3270 0.0700 ;
         RECT 0.3250 0.0560 0.3470 0.0700 ;
         RECT 0.3250 0.0700 0.3470 0.1120 ;
        RECT 0.0330 0.0880 0.2400 0.1040 ;
  END
END NAND3_X2

MACRO NAND4_X1
  CLASS core ;
  FOREIGN NAND4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.2940 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.2410 0.1280 0.2630 0.2870 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1570 0.1210 0.1790 0.2560 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1150 0.0970 0.1370 0.2240 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.0970 0.0530 0.2870 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.2560 0.0950 0.3220 ;
         RECT 0.0730 0.3220 0.0950 0.3520 ;
        RECT 0.0930 0.3220 0.2010 0.3520 ;
         RECT 0.1990 0.0820 0.2210 0.0960 ;
         RECT 0.1990 0.0960 0.2210 0.2560 ;
         RECT 0.1990 0.2560 0.2210 0.3220 ;
         RECT 0.1990 0.3220 0.2210 0.3520 ;
         RECT 0.2185 0.0820 0.2405 0.0960 ;
        RECT 0.2400 0.0320 0.2640 0.0820 ;
        RECT 0.2400 0.0820 0.2640 0.0960 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.3010 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.3010 0.0140 ;
    END
  END VSS
END NAND4_X1

MACRO NAND4_X2
  CLASS core ;
  FOREIGN NAND4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.4620 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.3660 0.1790 0.3900 0.2560 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.2410 0.1700 0.2630 0.2630 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1150 0.1210 0.1370 0.2560 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1280 0.0530 0.2560 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.2780 0.0950 0.2880 ;
         RECT 0.0730 0.2880 0.0950 0.3190 ;
         RECT 0.0730 0.3190 0.0950 0.3330 ;
        RECT 0.0940 0.3190 0.2850 0.3330 ;
         RECT 0.2830 0.1470 0.3050 0.1610 ;
         RECT 0.2830 0.1610 0.3050 0.2740 ;
         RECT 0.2830 0.2740 0.3050 0.2780 ;
         RECT 0.2830 0.2780 0.3050 0.2880 ;
         RECT 0.2830 0.3190 0.3050 0.3330 ;
        RECT 0.3030 0.1470 0.3690 0.1610 ;
        RECT 0.3030 0.2740 0.3690 0.2780 ;
        RECT 0.3030 0.2780 0.3690 0.2880 ;
        RECT 0.3030 0.3190 0.3690 0.3330 ;
         RECT 0.3670 0.1470 0.3890 0.1610 ;
         RECT 0.3670 0.2740 0.3890 0.2780 ;
         RECT 0.3670 0.2780 0.3890 0.2880 ;
         RECT 0.3670 0.2880 0.3890 0.3190 ;
         RECT 0.3670 0.3190 0.3890 0.3330 ;
        RECT 0.3870 0.1470 0.4290 0.1610 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.4300 0.3980 ;
        RECT 0.4300 0.3700 0.4690 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.4690 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0310 0.0510 0.0530 0.0650 ;
         RECT 0.0310 0.0650 0.0530 0.1060 ;
        RECT 0.0520 0.0510 0.2820 0.0650 ;
        RECT 0.1800 0.1150 0.4090 0.1290 ;
         RECT 0.4085 0.0320 0.4305 0.1150 ;
         RECT 0.4085 0.1150 0.4305 0.1290 ;
        RECT 0.0960 0.0830 0.3240 0.0970 ;
      LAYER M1 ;
         RECT 0.0310 0.0510 0.0530 0.0650 ;
         RECT 0.0310 0.0650 0.0530 0.1060 ;
        RECT 0.0520 0.0510 0.2820 0.0650 ;
        RECT 0.1800 0.1150 0.4090 0.1290 ;
         RECT 0.4085 0.0320 0.4305 0.1150 ;
         RECT 0.4085 0.1150 0.4305 0.1290 ;
        RECT 0.0960 0.0830 0.3240 0.0970 ;
  END
END NAND4_X2

MACRO NOR2_X1
  CLASS core ;
  FOREIGN NOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.1680 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1150 0.0970 0.1370 0.2560 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.0970 0.0530 0.2560 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.0650 0.0950 0.2880 ;
         RECT 0.0730 0.2880 0.0950 0.3180 ;
        RECT 0.0930 0.2880 0.1150 0.3180 ;
         RECT 0.1145 0.2880 0.1365 0.3180 ;
         RECT 0.1145 0.3180 0.1365 0.3520 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.1750 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.1750 0.0140 ;
    END
  END VSS
END NOR2_X1

MACRO NOR2_X2
  CLASS core ;
  FOREIGN NOR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.2520 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1150 0.1080 0.1370 0.2560 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.0320 0.0530 0.0460 ;
         RECT 0.0310 0.0460 0.0530 0.2470 ;
        RECT 0.0510 0.0320 0.2010 0.0460 ;
         RECT 0.1990 0.0320 0.2210 0.0460 ;
         RECT 0.1990 0.0460 0.2210 0.2470 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.0640 0.0950 0.0780 ;
         RECT 0.0730 0.0780 0.0950 0.1720 ;
         RECT 0.0730 0.1720 0.0950 0.2780 ;
         RECT 0.0730 0.2780 0.0950 0.2920 ;
        RECT 0.0930 0.0640 0.1150 0.0780 ;
        RECT 0.0930 0.2780 0.1150 0.2920 ;
         RECT 0.1145 0.0640 0.1365 0.0780 ;
         RECT 0.1145 0.2780 0.1365 0.2920 ;
         RECT 0.1145 0.2920 0.1365 0.3200 ;
        RECT 0.1360 0.0640 0.1590 0.0780 ;
         RECT 0.1570 0.0640 0.1790 0.0780 ;
         RECT 0.1570 0.0780 0.1790 0.1720 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.2590 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.2590 0.0140 ;
    END
  END VSS
END NOR2_X2

MACRO NOR3_X1
  CLASS core ;
  FOREIGN NOR3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.2520 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1570 0.1600 0.1790 0.2240 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1150 0.0970 0.1370 0.2760 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.0970 0.0530 0.2760 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.0320 0.0950 0.0460 ;
         RECT 0.0730 0.0460 0.0950 0.1280 ;
         RECT 0.0730 0.1280 0.0950 0.2560 ;
         RECT 0.0730 0.2560 0.0950 0.3070 ;
         RECT 0.0730 0.3070 0.0950 0.3210 ;
        RECT 0.0930 0.0320 0.1990 0.0460 ;
        RECT 0.0930 0.3070 0.1990 0.3210 ;
         RECT 0.1985 0.0320 0.2205 0.0460 ;
         RECT 0.1985 0.0460 0.2205 0.1280 ;
         RECT 0.1985 0.2560 0.2205 0.3070 ;
         RECT 0.1985 0.3070 0.2205 0.3210 ;
         RECT 0.1985 0.3210 0.2205 0.3520 ;
         RECT 0.2095 0.0320 0.2315 0.0460 ;
         RECT 0.2095 0.0460 0.2315 0.1280 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.2590 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.2590 0.0140 ;
    END
  END VSS
END NOR3_X1

MACRO NOR3_X2
  CLASS core ;
  FOREIGN NOR3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.3780 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.3250 0.1280 0.3470 0.2240 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1990 0.1280 0.2210 0.2560 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1280 0.0530 0.2600 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.0560 0.0770 0.2850 0.1060 ;
         RECT 0.2830 0.0770 0.3050 0.1060 ;
         RECT 0.2830 0.1060 0.3050 0.2880 ;
         RECT 0.3015 0.0770 0.3235 0.1060 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.3450 0.3980 ;
        RECT 0.3450 0.3700 0.3850 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.3850 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.1380 0.3140 0.3270 0.3280 ;
         RECT 0.3250 0.2580 0.3470 0.3140 ;
         RECT 0.3250 0.3140 0.3470 0.3280 ;
        RECT 0.0560 0.2780 0.2490 0.2960 ;
      LAYER M1 ;
        RECT 0.1380 0.3140 0.3270 0.3280 ;
         RECT 0.3250 0.2580 0.3470 0.3140 ;
         RECT 0.3250 0.3140 0.3470 0.3280 ;
        RECT 0.0560 0.2780 0.2490 0.2960 ;
  END
END NOR3_X2

MACRO NOR4_X1
  CLASS core ;
  FOREIGN NOR4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.2940 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.2410 0.0970 0.2630 0.2560 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1570 0.0970 0.1790 0.2560 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1150 0.1280 0.1370 0.2870 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.0970 0.0530 0.2870 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.0320 0.0950 0.0510 ;
         RECT 0.0730 0.0510 0.0950 0.1080 ;
        RECT 0.0930 0.0320 0.2010 0.0510 ;
         RECT 0.1990 0.0320 0.2210 0.0510 ;
         RECT 0.1990 0.0510 0.2210 0.1080 ;
         RECT 0.1990 0.1080 0.2210 0.2880 ;
         RECT 0.1990 0.2880 0.2210 0.3020 ;
         RECT 0.2185 0.2880 0.2405 0.3020 ;
        RECT 0.2400 0.2880 0.2640 0.3020 ;
        RECT 0.2400 0.3020 0.2640 0.3520 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.3010 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.3010 0.0140 ;
    END
  END VSS
END NOR4_X1

MACRO NOR4_X2
  CLASS core ;
  FOREIGN NOR4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.4620 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.3660 0.1280 0.3900 0.2030 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.2410 0.1210 0.2630 0.2190 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1570 0.1210 0.1790 0.2630 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1150 0.1280 0.1370 0.2580 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.0510 0.0950 0.0650 ;
         RECT 0.0730 0.0650 0.0950 0.0960 ;
         RECT 0.0730 0.0960 0.0950 0.1060 ;
        RECT 0.0940 0.0510 0.2850 0.0650 ;
         RECT 0.2830 0.0510 0.3050 0.0650 ;
         RECT 0.2830 0.0960 0.3050 0.1060 ;
         RECT 0.2830 0.1060 0.3050 0.1100 ;
         RECT 0.2830 0.1100 0.3050 0.2210 ;
         RECT 0.2830 0.2210 0.3050 0.2350 ;
        RECT 0.3030 0.0510 0.3690 0.0650 ;
        RECT 0.3030 0.0960 0.3690 0.1060 ;
        RECT 0.3030 0.1060 0.3690 0.1100 ;
        RECT 0.3030 0.2210 0.3690 0.2350 ;
         RECT 0.3670 0.0510 0.3890 0.0650 ;
         RECT 0.3670 0.0650 0.3890 0.0960 ;
         RECT 0.3670 0.0960 0.3890 0.1060 ;
         RECT 0.3670 0.1060 0.3890 0.1100 ;
         RECT 0.3670 0.2210 0.3890 0.2350 ;
        RECT 0.3870 0.2210 0.4350 0.2350 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.2820 0.3980 ;
        RECT 0.2820 0.3700 0.3240 0.3980 ;
        RECT 0.3240 0.3700 0.4300 0.3980 ;
        RECT 0.4300 0.3700 0.4690 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.4690 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.1380 0.2850 0.3240 0.3010 ;
         RECT 0.0310 0.2780 0.0530 0.3190 ;
         RECT 0.0310 0.3190 0.0530 0.3330 ;
        RECT 0.0520 0.3190 0.2820 0.3330 ;
        RECT 0.2220 0.2530 0.4090 0.2670 ;
         RECT 0.4085 0.2530 0.4305 0.2670 ;
         RECT 0.4085 0.2670 0.4305 0.3430 ;
      LAYER M1 ;
        RECT 0.1380 0.2850 0.3240 0.3010 ;
         RECT 0.0310 0.2780 0.0530 0.3190 ;
         RECT 0.0310 0.3190 0.0530 0.3330 ;
        RECT 0.0520 0.3190 0.2820 0.3330 ;
        RECT 0.2220 0.2530 0.4090 0.2670 ;
         RECT 0.4085 0.2530 0.4305 0.2670 ;
         RECT 0.4085 0.2670 0.4305 0.3430 ;
  END
END NOR4_X2

MACRO OAI21_X1
  CLASS core ;
  FOREIGN OAI21_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.2520 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1150 0.1280 0.1370 0.2880 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1280 0.0530 0.3170 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1990 0.1280 0.2210 0.2880 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.1280 0.0950 0.3180 ;
         RECT 0.0730 0.3180 0.0950 0.3340 ;
        RECT 0.0930 0.3180 0.1960 0.3340 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.1960 0.3980 ;
        RECT 0.1960 0.3700 0.2590 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.2590 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0310 0.0360 0.0530 0.0780 ;
         RECT 0.0310 0.0780 0.0530 0.0940 ;
        RECT 0.0510 0.0780 0.1960 0.0940 ;
      LAYER M1 ;
         RECT 0.0310 0.0360 0.0530 0.0780 ;
         RECT 0.0310 0.0780 0.0530 0.0940 ;
        RECT 0.0510 0.0780 0.1960 0.0940 ;
  END
END OAI21_X1

MACRO OAI21_X2
  CLASS core ;
  FOREIGN OAI21_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.3780 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.2400 0.1600 0.2640 0.2240 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1570 0.1210 0.1790 0.1410 ;
         RECT 0.1570 0.1410 0.1790 0.2510 ;
         RECT 0.1570 0.2510 0.1790 0.2650 ;
        RECT 0.1770 0.2510 0.3270 0.2650 ;
         RECT 0.3250 0.1410 0.3470 0.2510 ;
         RECT 0.3250 0.2510 0.3470 0.2650 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.1280 0.0950 0.2620 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.0190 0.2850 0.1170 0.3010 ;
         RECT 0.1150 0.0830 0.1370 0.0970 ;
         RECT 0.1150 0.0970 0.1370 0.1390 ;
         RECT 0.1150 0.1390 0.1370 0.2850 ;
         RECT 0.1150 0.2850 0.1370 0.3010 ;
        RECT 0.1350 0.0830 0.2800 0.0970 ;
        RECT 0.1350 0.2850 0.2800 0.3010 ;
         RECT 0.2715 0.0830 0.2935 0.0970 ;
         RECT 0.2830 0.0830 0.3050 0.0970 ;
         RECT 0.2830 0.0970 0.3050 0.1390 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.3510 0.3980 ;
        RECT 0.3510 0.3700 0.3850 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.3850 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0310 0.0510 0.0530 0.0650 ;
         RECT 0.0310 0.0650 0.0530 0.1060 ;
        RECT 0.0520 0.0510 0.3270 0.0650 ;
         RECT 0.3250 0.0510 0.3470 0.0650 ;
         RECT 0.3250 0.0650 0.3470 0.1060 ;
         RECT 0.3250 0.1060 0.3470 0.1080 ;
        RECT 0.0960 0.3190 0.3510 0.3330 ;
      LAYER M1 ;
         RECT 0.0310 0.0510 0.0530 0.0650 ;
         RECT 0.0310 0.0650 0.0530 0.1060 ;
        RECT 0.0520 0.0510 0.3270 0.0650 ;
         RECT 0.3250 0.0510 0.3470 0.0650 ;
         RECT 0.3250 0.0650 0.3470 0.1060 ;
         RECT 0.3250 0.1060 0.3470 0.1080 ;
        RECT 0.0960 0.3190 0.3510 0.3330 ;
  END
END OAI21_X2

MACRO OAI22_X1
  CLASS core ;
  FOREIGN OAI22_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.2940 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1570 0.1000 0.1790 0.2880 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.2410 0.1400 0.2630 0.2880 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1150 0.0960 0.1370 0.2560 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.0960 0.0530 0.2880 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.0920 0.3190 0.2010 0.3330 ;
         RECT 0.1990 0.0910 0.2210 0.3190 ;
         RECT 0.1990 0.3190 0.2210 0.3330 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.2610 0.3980 ;
        RECT 0.2610 0.3700 0.3010 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.3010 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.0330 0.0500 0.2430 0.0660 ;
         RECT 0.2410 0.0500 0.2630 0.0660 ;
         RECT 0.2410 0.0660 0.2630 0.1060 ;
      LAYER M1 ;
        RECT 0.0330 0.0500 0.2430 0.0660 ;
         RECT 0.2410 0.0500 0.2630 0.0660 ;
         RECT 0.2410 0.0660 0.2630 0.1060 ;
  END
END OAI22_X1

MACRO OAI22_X2
  CLASS core ;
  FOREIGN OAI22_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.5040 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.2830 0.1280 0.3050 0.1400 ;
         RECT 0.2830 0.1400 0.3050 0.2330 ;
         RECT 0.2830 0.2330 0.3050 0.2470 ;
        RECT 0.3030 0.2330 0.4530 0.2470 ;
         RECT 0.4510 0.1400 0.4730 0.2330 ;
         RECT 0.4510 0.2330 0.4730 0.2470 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.3670 0.1280 0.3890 0.1990 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1990 0.1210 0.2210 0.2430 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.1210 0.0950 0.2560 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1570 0.1930 0.1790 0.2650 ;
         RECT 0.1570 0.2650 0.1790 0.2790 ;
        RECT 0.1770 0.2650 0.2430 0.2790 ;
         RECT 0.2410 0.0840 0.2630 0.0980 ;
         RECT 0.2410 0.0980 0.2630 0.1390 ;
         RECT 0.2410 0.1390 0.2630 0.1930 ;
         RECT 0.2410 0.1930 0.2630 0.2650 ;
         RECT 0.2410 0.2650 0.2630 0.2790 ;
        RECT 0.2610 0.0840 0.4110 0.0980 ;
        RECT 0.2610 0.2650 0.4110 0.2790 ;
         RECT 0.4090 0.0840 0.4310 0.0980 ;
         RECT 0.4090 0.0980 0.4310 0.1390 ;
         RECT 0.4090 0.2650 0.4310 0.2790 ;
        RECT 0.4290 0.2650 0.4530 0.2790 ;
         RECT 0.4510 0.2650 0.4730 0.2790 ;
         RECT 0.4510 0.2790 0.4730 0.3360 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.2380 0.3980 ;
        RECT 0.2380 0.3700 0.4290 0.3980 ;
        RECT 0.4290 0.3700 0.4710 0.3980 ;
        RECT 0.4710 0.3700 0.5110 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.5110 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.2640 0.3020 0.4110 0.3180 ;
         RECT 0.4090 0.3020 0.4310 0.3180 ;
         RECT 0.4090 0.3180 0.4310 0.3480 ;
        RECT 0.0270 0.0500 0.4530 0.0660 ;
         RECT 0.4510 0.0500 0.4730 0.0660 ;
         RECT 0.4510 0.0660 0.4730 0.1060 ;
        RECT 0.0330 0.3060 0.2380 0.3350 ;
      LAYER M1 ;
        RECT 0.2640 0.3020 0.4110 0.3180 ;
         RECT 0.4090 0.3020 0.4310 0.3180 ;
         RECT 0.4090 0.3180 0.4310 0.3480 ;
        RECT 0.0270 0.0500 0.4530 0.0660 ;
         RECT 0.4510 0.0500 0.4730 0.0660 ;
         RECT 0.4510 0.0660 0.4730 0.1060 ;
        RECT 0.0330 0.3060 0.2380 0.3350 ;
  END
END OAI22_X2

MACRO OR2_X1
  CLASS core ;
  FOREIGN OR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.2520 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1150 0.0480 0.1370 0.2560 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1220 0.0530 0.3200 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1990 0.0570 0.2210 0.3200 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.1770 0.3980 ;
        RECT 0.1770 0.3700 0.2590 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.2590 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0730 0.0650 0.0950 0.1680 ;
         RECT 0.0730 0.1680 0.0950 0.2780 ;
         RECT 0.0730 0.2780 0.0950 0.2920 ;
        RECT 0.0930 0.2780 0.1590 0.2920 ;
         RECT 0.1570 0.1680 0.1790 0.2780 ;
         RECT 0.1570 0.2780 0.1790 0.2920 ;
      LAYER M1 ;
         RECT 0.0730 0.0650 0.0950 0.1680 ;
         RECT 0.0730 0.1680 0.0950 0.2780 ;
         RECT 0.0730 0.2780 0.0950 0.2920 ;
        RECT 0.0930 0.2780 0.1590 0.2920 ;
         RECT 0.1570 0.1680 0.1790 0.2780 ;
         RECT 0.1570 0.2780 0.1790 0.2920 ;
  END
END OR2_X1

MACRO OR2_X2
  CLASS core ;
  FOREIGN OR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.2940 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.1210 0.0950 0.2560 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1280 0.0530 0.2560 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1885 0.0320 0.2105 0.0680 ;
         RECT 0.1885 0.3190 0.2105 0.3520 ;
         RECT 0.1990 0.0320 0.2210 0.0680 ;
         RECT 0.1990 0.0680 0.2210 0.3190 ;
         RECT 0.1990 0.3190 0.2210 0.3520 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.1770 0.3980 ;
        RECT 0.1770 0.3700 0.3010 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.3010 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.0510 0.0770 0.0960 0.0940 ;
        RECT 0.0960 0.0770 0.1590 0.0940 ;
        RECT 0.0960 0.2900 0.1590 0.3040 ;
         RECT 0.1570 0.0770 0.1790 0.0940 ;
         RECT 0.1570 0.0940 0.1790 0.2900 ;
         RECT 0.1570 0.2900 0.1790 0.3040 ;
      LAYER M1 ;
        RECT 0.0510 0.0770 0.0960 0.0940 ;
        RECT 0.0960 0.0770 0.1590 0.0940 ;
        RECT 0.0960 0.2900 0.1590 0.3040 ;
         RECT 0.1570 0.0770 0.1790 0.0940 ;
         RECT 0.1570 0.0940 0.1790 0.2900 ;
         RECT 0.1570 0.2900 0.1790 0.3040 ;
  END
END OR2_X2

MACRO OR3_X1
  CLASS core ;
  FOREIGN OR3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.3360 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1990 0.0960 0.2210 0.2880 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1145 0.0960 0.1365 0.2880 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.0300 0.0960 0.0540 0.2880 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.2830 0.0570 0.3050 0.3270 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.1540 0.3980 ;
        RECT 0.1540 0.3700 0.2610 0.3980 ;
        RECT 0.2610 0.3700 0.3430 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.3430 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.0350 0.0540 0.1820 0.0680 ;
        RECT 0.1820 0.0540 0.2430 0.0680 ;
        RECT 0.1820 0.3160 0.2430 0.3360 ;
         RECT 0.2410 0.0540 0.2630 0.0680 ;
         RECT 0.2410 0.0680 0.2630 0.3160 ;
         RECT 0.2410 0.3160 0.2630 0.3360 ;
        RECT 0.0560 0.3180 0.1540 0.3340 ;
      LAYER M1 ;
        RECT 0.0350 0.0540 0.1820 0.0680 ;
        RECT 0.1820 0.0540 0.2430 0.0680 ;
        RECT 0.1820 0.3160 0.2430 0.3360 ;
         RECT 0.2410 0.0540 0.2630 0.0680 ;
         RECT 0.2410 0.0680 0.2630 0.3160 ;
         RECT 0.2410 0.3160 0.2630 0.3360 ;
        RECT 0.0560 0.3180 0.1540 0.3340 ;
  END
END OR3_X1

MACRO OR3_X2
  CLASS core ;
  FOREIGN OR3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.3360 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.1280 0.0950 0.2240 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1280 0.0530 0.2630 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1570 0.1160 0.1790 0.2240 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.2305 0.0320 0.2525 0.0650 ;
         RECT 0.2305 0.3180 0.2525 0.3520 ;
         RECT 0.2410 0.0320 0.2630 0.0650 ;
         RECT 0.2410 0.0650 0.2630 0.3180 ;
         RECT 0.2410 0.3180 0.2630 0.3520 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.1980 0.3980 ;
         RECT 0.1975 0.3700 0.2195 0.3980 ;
        RECT 0.2190 0.3700 0.3430 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.3430 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0310 0.2860 0.0530 0.3020 ;
         RECT 0.0310 0.3020 0.0530 0.3430 ;
        RECT 0.0510 0.2860 0.1980 0.3020 ;
        RECT 0.0390 0.0780 0.0920 0.0940 ;
        RECT 0.0920 0.0780 0.2010 0.0940 ;
        RECT 0.0920 0.2520 0.2010 0.2680 ;
         RECT 0.1990 0.0780 0.2210 0.0940 ;
         RECT 0.1990 0.0940 0.2210 0.2520 ;
         RECT 0.1990 0.2520 0.2210 0.2680 ;
      LAYER M1 ;
         RECT 0.0310 0.2860 0.0530 0.3020 ;
         RECT 0.0310 0.3020 0.0530 0.3430 ;
        RECT 0.0510 0.2860 0.1980 0.3020 ;
        RECT 0.0390 0.0780 0.0920 0.0940 ;
        RECT 0.0920 0.0780 0.2010 0.0940 ;
        RECT 0.0920 0.2520 0.2010 0.2680 ;
         RECT 0.1990 0.0780 0.2210 0.0940 ;
         RECT 0.1990 0.0940 0.2210 0.2520 ;
         RECT 0.1990 0.2520 0.2210 0.2680 ;
  END
END OR3_X2

MACRO OR4_X1
  CLASS core ;
  FOREIGN OR4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.3780 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.2410 0.0960 0.2630 0.2880 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1575 0.0960 0.1795 0.2880 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.0990 0.0950 0.2880 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.0960 0.0530 0.2880 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.3250 0.0570 0.3470 0.3200 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.1960 0.3980 ;
        RECT 0.1960 0.3700 0.3030 0.3980 ;
        RECT 0.3030 0.3700 0.3850 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.3850 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.0350 0.0510 0.2220 0.0650 ;
        RECT 0.2220 0.0510 0.2850 0.0650 ;
        RECT 0.2220 0.3150 0.2850 0.3310 ;
         RECT 0.2830 0.0510 0.3050 0.0650 ;
         RECT 0.2830 0.0650 0.3050 0.3150 ;
         RECT 0.2830 0.3150 0.3050 0.3310 ;
        RECT 0.0960 0.3080 0.1960 0.3280 ;
      LAYER M1 ;
        RECT 0.0350 0.0510 0.2220 0.0650 ;
        RECT 0.2220 0.0510 0.2850 0.0650 ;
        RECT 0.2220 0.3150 0.2850 0.3310 ;
         RECT 0.2830 0.0510 0.3050 0.0650 ;
         RECT 0.2830 0.0650 0.3050 0.3150 ;
         RECT 0.2830 0.3150 0.3050 0.3310 ;
        RECT 0.0960 0.3080 0.1960 0.3280 ;
  END
END OR4_X1

MACRO OR4_X2
  CLASS core ;
  FOREIGN OR4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.4200 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1990 0.0960 0.2210 0.2650 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1570 0.1060 0.1790 0.2880 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.1060 0.0950 0.2880 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.0960 0.0530 0.2880 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.3250 0.0640 0.3470 0.3520 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.1980 0.3980 ;
        RECT 0.1980 0.3700 0.3020 0.3980 ;
        RECT 0.3020 0.3700 0.4270 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.4270 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.0960 0.3120 0.1980 0.3400 ;
        RECT 0.0350 0.0430 0.2240 0.0720 ;
        RECT 0.2240 0.0430 0.2830 0.0720 ;
        RECT 0.2240 0.2840 0.2830 0.3120 ;
         RECT 0.2815 0.0430 0.3035 0.0720 ;
         RECT 0.2815 0.0720 0.3035 0.2840 ;
         RECT 0.2815 0.2840 0.3035 0.3120 ;
      LAYER M1 ;
        RECT 0.0960 0.3120 0.1980 0.3400 ;
        RECT 0.0350 0.0430 0.2240 0.0720 ;
        RECT 0.2240 0.0430 0.2830 0.0720 ;
        RECT 0.2240 0.2840 0.2830 0.3120 ;
         RECT 0.2815 0.0430 0.3035 0.0720 ;
         RECT 0.2815 0.0720 0.3035 0.2840 ;
         RECT 0.2815 0.2840 0.3035 0.3120 ;
  END
END OR4_X2

MACRO SDFFRNQ_X1
  CLASS core ;
  FOREIGN SDFFRNQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 1.2600 BY 0.3840 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.3215 0.1820 0.3435 0.2640 ;
         RECT 0.3305 0.1820 0.3525 0.2640 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
         RECT 0.6330 0.1640 0.9540 0.1880 ;
         RECT 0.9540 0.1640 1.0450 0.1880 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1990 0.1860 0.2210 0.2860 ;
         RECT 0.1990 0.2860 0.2210 0.3000 ;
        RECT 0.2190 0.2860 0.3380 0.3000 ;
        RECT 0.3380 0.2860 0.3690 0.3000 ;
         RECT 0.3670 0.1570 0.3890 0.1860 ;
         RECT 0.3670 0.1860 0.3890 0.2860 ;
         RECT 0.3670 0.2860 0.3890 0.3000 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.2410 0.1820 0.2630 0.2560 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1380 0.0530 0.2670 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 1.2075 0.0320 1.2295 0.3520 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.0930 0.3980 ;
        RECT 0.0930 0.3700 0.1350 0.3980 ;
        RECT 0.1350 0.3700 0.4950 0.3980 ;
         RECT 0.4930 0.3700 0.5150 0.3980 ;
        RECT 0.5130 0.3700 0.7000 0.3980 ;
        RECT 0.7000 0.3700 0.9330 0.3980 ;
        RECT 0.9330 0.3700 0.9780 0.3980 ;
        RECT 0.9780 0.3700 1.1430 0.3980 ;
        RECT 1.1430 0.3700 1.2670 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 1.2670 0.0140 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
         RECT 0.0960 0.2600 0.8700 0.2840 ;
         RECT 0.4740 0.1960 0.7360 0.2200 ;
         RECT 0.0540 0.1320 0.9540 0.1560 ;
      LAYER MINT1 ;
         RECT 0.0960 0.2600 0.8700 0.2840 ;
         RECT 0.4740 0.1960 0.7360 0.2200 ;
         RECT 0.0540 0.1320 0.9540 0.1560 ;
      LAYER M1 ;
        RECT 0.0300 0.0480 0.0540 0.1020 ;
        RECT 0.0300 0.1020 0.0540 0.1160 ;
        RECT 0.0300 0.3020 0.0540 0.3160 ;
        RECT 0.0300 0.3160 0.0540 0.3440 ;
         RECT 0.0535 0.1020 0.0755 0.1160 ;
         RECT 0.0535 0.3020 0.0755 0.3160 ;
         RECT 0.0730 0.1020 0.0950 0.1160 ;
         RECT 0.0730 0.1160 0.0950 0.3020 ;
         RECT 0.0730 0.3020 0.0950 0.3160 ;
         RECT 0.1570 0.0480 0.1790 0.1340 ;
         RECT 0.1570 0.1340 0.1790 0.1480 ;
         RECT 0.1570 0.1480 0.1790 0.3360 ;
        RECT 0.1770 0.1340 0.3380 0.1480 ;
        RECT 0.2220 0.0920 0.4110 0.1060 ;
         RECT 0.4090 0.0920 0.4310 0.1060 ;
         RECT 0.4090 0.1060 0.4310 0.1380 ;
        RECT 0.2570 0.3180 0.4950 0.3340 ;
         RECT 0.4930 0.1240 0.5150 0.2730 ;
        RECT 0.3060 0.0510 0.5760 0.0650 ;
        RECT 0.6960 0.1200 0.7210 0.2230 ;
         RECT 0.7870 0.0860 0.8090 0.2560 ;
         RECT 0.9565 0.0730 0.9785 0.3490 ;
        RECT 0.7650 0.3090 0.8730 0.3230 ;
         RECT 0.8710 0.0320 0.8930 0.0460 ;
         RECT 0.8710 0.0460 0.8930 0.1830 ;
         RECT 0.8710 0.1830 0.8930 0.3090 ;
         RECT 0.8710 0.3090 0.8930 0.3230 ;
        RECT 0.8910 0.0320 1.0550 0.0460 ;
         RECT 1.0530 0.0320 1.0750 0.0460 ;
         RECT 1.0530 0.0460 1.0750 0.1830 ;
         RECT 1.0180 0.2300 1.0400 0.3120 ;
         RECT 1.0180 0.3120 1.0400 0.3400 ;
        RECT 1.0380 0.3120 1.1250 0.3400 ;
         RECT 1.1230 0.0360 1.1450 0.2300 ;
         RECT 1.1230 0.2300 1.1450 0.3120 ;
         RECT 1.1230 0.3120 1.1450 0.3400 ;
         RECT 0.1150 0.0620 0.1370 0.2870 ;
         RECT 0.4510 0.1940 0.4730 0.2950 ;
         RECT 0.5365 0.1280 0.5585 0.2340 ;
         RECT 0.4510 0.0830 0.4730 0.0970 ;
         RECT 0.4510 0.0970 0.4730 0.1380 ;
        RECT 0.4710 0.0830 0.6180 0.0970 ;
        RECT 0.6500 0.1210 0.6730 0.2110 ;
        RECT 0.5180 0.3180 0.7000 0.3340 ;
         RECT 0.5915 0.1370 0.6135 0.2450 ;
         RECT 0.5915 0.2450 0.6135 0.2590 ;
        RECT 0.6120 0.2450 0.7440 0.2590 ;
         RECT 0.7435 0.0410 0.7655 0.1370 ;
         RECT 0.7435 0.1370 0.7655 0.2450 ;
         RECT 0.7435 0.2450 0.7655 0.2590 ;
         RECT 0.8290 0.0890 0.8510 0.2870 ;
         RECT 0.9130 0.0890 0.9350 0.2470 ;
        RECT 1.0050 0.0770 1.0310 0.2080 ;
      LAYER V1 ;
        RECT 0.0750 0.1370 0.0930 0.1510 ;
        RECT 0.1170 0.2650 0.1350 0.2790 ;
        RECT 0.4530 0.2650 0.4710 0.2790 ;
        RECT 0.4950 0.2010 0.5130 0.2150 ;
        RECT 0.5370 0.1370 0.5550 0.1510 ;
        RECT 0.6540 0.1690 0.6730 0.1830 ;
        RECT 0.6960 0.2010 0.7150 0.2150 ;
        RECT 0.7890 0.1370 0.8070 0.1510 ;
        RECT 0.8310 0.2650 0.8490 0.2790 ;
        RECT 0.9150 0.1370 0.9330 0.1510 ;
        RECT 1.0050 0.1690 1.0240 0.1830 ;
      LAYER M1 ;
        RECT 0.0300 0.0480 0.0540 0.1020 ;
        RECT 0.0300 0.1020 0.0540 0.1160 ;
        RECT 0.0300 0.3020 0.0540 0.3160 ;
        RECT 0.0300 0.3160 0.0540 0.3440 ;
         RECT 0.0535 0.1020 0.0755 0.1160 ;
         RECT 0.0535 0.3020 0.0755 0.3160 ;
         RECT 0.0730 0.1020 0.0950 0.1160 ;
         RECT 0.0730 0.1160 0.0950 0.3020 ;
         RECT 0.0730 0.3020 0.0950 0.3160 ;
         RECT 0.1570 0.0480 0.1790 0.1340 ;
         RECT 0.1570 0.1340 0.1790 0.1480 ;
         RECT 0.1570 0.1480 0.1790 0.3360 ;
        RECT 0.1770 0.1340 0.3380 0.1480 ;
        RECT 0.2220 0.0920 0.4110 0.1060 ;
         RECT 0.4090 0.0920 0.4310 0.1060 ;
         RECT 0.4090 0.1060 0.4310 0.1380 ;
        RECT 0.2570 0.3180 0.4950 0.3340 ;
         RECT 0.4930 0.1240 0.5150 0.2730 ;
        RECT 0.3060 0.0510 0.5760 0.0650 ;
        RECT 0.6960 0.1200 0.7210 0.2230 ;
         RECT 0.7870 0.0860 0.8090 0.2560 ;
         RECT 0.9565 0.0730 0.9785 0.3490 ;
        RECT 0.7650 0.3090 0.8730 0.3230 ;
         RECT 0.8710 0.0320 0.8930 0.0460 ;
         RECT 0.8710 0.0460 0.8930 0.1830 ;
         RECT 0.8710 0.1830 0.8930 0.3090 ;
         RECT 0.8710 0.3090 0.8930 0.3230 ;
        RECT 0.8910 0.0320 1.0550 0.0460 ;
         RECT 1.0530 0.0320 1.0750 0.0460 ;
         RECT 1.0530 0.0460 1.0750 0.1830 ;
         RECT 1.0180 0.2300 1.0400 0.3120 ;
         RECT 1.0180 0.3120 1.0400 0.3400 ;
        RECT 1.0380 0.3120 1.1250 0.3400 ;
         RECT 1.1230 0.0360 1.1450 0.2300 ;
         RECT 1.1230 0.2300 1.1450 0.3120 ;
         RECT 1.1230 0.3120 1.1450 0.3400 ;
         RECT 0.1150 0.0620 0.1370 0.2870 ;
         RECT 0.4510 0.1940 0.4730 0.2950 ;
         RECT 0.5365 0.1280 0.5585 0.2340 ;
         RECT 0.4510 0.0830 0.4730 0.0970 ;
         RECT 0.4510 0.0970 0.4730 0.1380 ;
        RECT 0.4710 0.0830 0.6180 0.0970 ;
        RECT 0.6500 0.1210 0.6730 0.2110 ;
        RECT 0.5180 0.3180 0.7000 0.3340 ;
         RECT 0.5915 0.1370 0.6135 0.2450 ;
         RECT 0.5915 0.2450 0.6135 0.2590 ;
        RECT 0.6120 0.2450 0.7440 0.2590 ;
         RECT 0.7435 0.0410 0.7655 0.1370 ;
         RECT 0.7435 0.1370 0.7655 0.2450 ;
         RECT 0.7435 0.2450 0.7655 0.2590 ;
         RECT 0.8290 0.0890 0.8510 0.2870 ;
         RECT 0.9130 0.0890 0.9350 0.2470 ;
        RECT 1.0050 0.0770 1.0310 0.2080 ;
  END
END SDFFRNQ_X1

MACRO SDFFSNQ_X1
  CLASS core ;
  FOREIGN SDFFSNQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 1.2600 BY 0.3840 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.3200 0.1920 0.3420 0.2640 ;
         RECT 0.3290 0.1920 0.3510 0.2640 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1990 0.1860 0.2210 0.2860 ;
         RECT 0.1990 0.2860 0.2210 0.3000 ;
        RECT 0.2190 0.2860 0.3350 0.3000 ;
        RECT 0.3350 0.2860 0.3690 0.3000 ;
         RECT 0.3670 0.1570 0.3890 0.1860 ;
         RECT 0.3670 0.1860 0.3890 0.2860 ;
         RECT 0.3670 0.2860 0.3890 0.3000 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.2410 0.1820 0.2630 0.2560 ;
    END
  END SI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
         RECT 0.6290 0.1640 0.9540 0.1880 ;
         RECT 0.9540 0.1640 1.0410 0.1880 ;
    END
  END SN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1360 0.0530 0.2560 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 1.2075 0.0320 1.2295 0.3520 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.0930 0.3980 ;
        RECT 0.0930 0.3700 0.1350 0.3980 ;
        RECT 0.1350 0.3700 0.4900 0.3980 ;
        RECT 0.4900 0.3700 0.5130 0.3980 ;
        RECT 0.5130 0.3700 0.5660 0.3980 ;
        RECT 0.5660 0.3700 1.0800 0.3980 ;
        RECT 1.0800 0.3700 1.1430 0.3980 ;
        RECT 1.1430 0.3700 1.2670 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 1.2670 0.0140 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
         RECT 0.0960 0.2600 0.8700 0.2840 ;
         RECT 0.4740 0.1960 0.7310 0.2200 ;
         RECT 0.0540 0.1320 0.9540 0.1560 ;
      LAYER MINT1 ;
         RECT 0.0960 0.2600 0.8700 0.2840 ;
         RECT 0.4740 0.1960 0.7310 0.2200 ;
         RECT 0.0540 0.1320 0.9540 0.1560 ;
      LAYER M1 ;
         RECT 0.0310 0.0320 0.0530 0.1000 ;
         RECT 0.0310 0.1000 0.0530 0.1140 ;
         RECT 0.0310 0.3020 0.0530 0.3160 ;
         RECT 0.0310 0.3160 0.0530 0.3440 ;
        RECT 0.0520 0.1000 0.0750 0.1140 ;
        RECT 0.0520 0.3020 0.0750 0.3160 ;
         RECT 0.0730 0.1000 0.0950 0.1140 ;
         RECT 0.0730 0.1140 0.0950 0.3020 ;
         RECT 0.0730 0.3020 0.0950 0.3160 ;
         RECT 0.1570 0.0410 0.1790 0.1330 ;
         RECT 0.1570 0.1330 0.1790 0.1480 ;
         RECT 0.1570 0.1480 0.1790 0.3430 ;
        RECT 0.1770 0.1330 0.2850 0.1480 ;
        RECT 0.2850 0.1330 0.3350 0.1480 ;
        RECT 0.2220 0.0920 0.4110 0.1060 ;
         RECT 0.4090 0.0920 0.4310 0.1060 ;
         RECT 0.4090 0.1060 0.4310 0.1380 ;
        RECT 0.2570 0.3180 0.4900 0.3340 ;
         RECT 0.4930 0.1190 0.5150 0.2740 ;
        RECT 0.3060 0.0510 0.5760 0.0650 ;
        RECT 0.6430 0.1610 0.6680 0.2100 ;
         RECT 0.5875 0.1370 0.6095 0.2440 ;
         RECT 0.5875 0.2440 0.6095 0.2580 ;
        RECT 0.6080 0.2440 0.6620 0.2580 ;
         RECT 0.6610 0.2440 0.6830 0.2580 ;
         RECT 0.6610 0.2580 0.6830 0.3520 ;
        RECT 0.6820 0.2440 0.7470 0.2580 ;
         RECT 0.7450 0.0490 0.7670 0.1370 ;
         RECT 0.7450 0.1370 0.7670 0.2440 ;
         RECT 0.7450 0.2440 0.7670 0.2580 ;
         RECT 0.8290 0.0890 0.8510 0.2870 ;
         RECT 0.9130 0.0890 0.9350 0.2010 ;
         RECT 0.9995 0.0920 1.0215 0.2020 ;
        RECT 0.9200 0.3190 1.0800 0.3330 ;
         RECT 0.1150 0.0480 0.1370 0.3100 ;
         RECT 0.4275 0.1940 0.4495 0.2870 ;
         RECT 0.5445 0.1280 0.5665 0.2340 ;
         RECT 0.4510 0.0830 0.4730 0.0970 ;
         RECT 0.4510 0.0970 0.4730 0.1380 ;
        RECT 0.4710 0.0830 0.6180 0.0970 ;
        RECT 0.6920 0.1200 0.7170 0.2230 ;
         RECT 0.7870 0.0860 0.8090 0.1920 ;
        RECT 0.7650 0.3090 0.8730 0.3230 ;
         RECT 0.8710 0.0410 0.8930 0.0550 ;
         RECT 0.8710 0.0550 0.8930 0.1830 ;
         RECT 0.8710 0.1830 0.8930 0.3090 ;
         RECT 0.8710 0.3090 0.8930 0.3230 ;
        RECT 0.8910 0.0410 1.0550 0.0550 ;
        RECT 1.0550 0.0410 1.0800 0.0550 ;
        RECT 1.0550 0.0550 1.0800 0.1830 ;
         RECT 0.9575 0.2010 0.9795 0.2870 ;
         RECT 0.9575 0.2870 0.9795 0.3010 ;
        RECT 0.9780 0.2870 1.1250 0.3010 ;
         RECT 1.1230 0.0480 1.1450 0.2010 ;
         RECT 1.1230 0.2010 1.1450 0.2870 ;
         RECT 1.1230 0.2870 1.1450 0.3010 ;
      LAYER V1 ;
        RECT 0.0750 0.1370 0.0930 0.1510 ;
        RECT 0.1170 0.2650 0.1350 0.2790 ;
        RECT 0.4290 0.2650 0.4480 0.2790 ;
        RECT 0.4950 0.2010 0.5130 0.2150 ;
        RECT 0.5470 0.1370 0.5660 0.1510 ;
        RECT 0.6500 0.1690 0.6680 0.1830 ;
        RECT 0.6920 0.2010 0.7100 0.2150 ;
        RECT 0.7890 0.1370 0.8070 0.1510 ;
        RECT 0.8310 0.2650 0.8490 0.2790 ;
        RECT 0.9150 0.1370 0.9330 0.1510 ;
        RECT 1.0010 0.1690 1.0200 0.1830 ;
      LAYER M1 ;
         RECT 0.0310 0.0320 0.0530 0.1000 ;
         RECT 0.0310 0.1000 0.0530 0.1140 ;
         RECT 0.0310 0.3020 0.0530 0.3160 ;
         RECT 0.0310 0.3160 0.0530 0.3440 ;
        RECT 0.0520 0.1000 0.0750 0.1140 ;
        RECT 0.0520 0.3020 0.0750 0.3160 ;
         RECT 0.0730 0.1000 0.0950 0.1140 ;
         RECT 0.0730 0.1140 0.0950 0.3020 ;
         RECT 0.0730 0.3020 0.0950 0.3160 ;
         RECT 0.1570 0.0410 0.1790 0.1330 ;
         RECT 0.1570 0.1330 0.1790 0.1480 ;
         RECT 0.1570 0.1480 0.1790 0.3430 ;
        RECT 0.1770 0.1330 0.2850 0.1480 ;
        RECT 0.2850 0.1330 0.3350 0.1480 ;
        RECT 0.2220 0.0920 0.4110 0.1060 ;
         RECT 0.4090 0.0920 0.4310 0.1060 ;
         RECT 0.4090 0.1060 0.4310 0.1380 ;
        RECT 0.2570 0.3180 0.4900 0.3340 ;
         RECT 0.4930 0.1190 0.5150 0.2740 ;
        RECT 0.3060 0.0510 0.5760 0.0650 ;
        RECT 0.6430 0.1610 0.6680 0.2100 ;
         RECT 0.5875 0.1370 0.6095 0.2440 ;
         RECT 0.5875 0.2440 0.6095 0.2580 ;
        RECT 0.6080 0.2440 0.6620 0.2580 ;
         RECT 0.6610 0.2440 0.6830 0.2580 ;
         RECT 0.6610 0.2580 0.6830 0.3520 ;
        RECT 0.6820 0.2440 0.7470 0.2580 ;
         RECT 0.7450 0.0490 0.7670 0.1370 ;
         RECT 0.7450 0.1370 0.7670 0.2440 ;
         RECT 0.7450 0.2440 0.7670 0.2580 ;
         RECT 0.8290 0.0890 0.8510 0.2870 ;
         RECT 0.9130 0.0890 0.9350 0.2010 ;
         RECT 0.9995 0.0920 1.0215 0.2020 ;
        RECT 0.9200 0.3190 1.0800 0.3330 ;
         RECT 0.1150 0.0480 0.1370 0.3100 ;
         RECT 0.4275 0.1940 0.4495 0.2870 ;
         RECT 0.5445 0.1280 0.5665 0.2340 ;
         RECT 0.4510 0.0830 0.4730 0.0970 ;
         RECT 0.4510 0.0970 0.4730 0.1380 ;
        RECT 0.4710 0.0830 0.6180 0.0970 ;
        RECT 0.6920 0.1200 0.7170 0.2230 ;
         RECT 0.7870 0.0860 0.8090 0.1920 ;
        RECT 0.7650 0.3090 0.8730 0.3230 ;
         RECT 0.8710 0.0410 0.8930 0.0550 ;
         RECT 0.8710 0.0550 0.8930 0.1830 ;
         RECT 0.8710 0.1830 0.8930 0.3090 ;
         RECT 0.8710 0.3090 0.8930 0.3230 ;
        RECT 0.8910 0.0410 1.0550 0.0550 ;
        RECT 1.0550 0.0410 1.0800 0.0550 ;
        RECT 1.0550 0.0550 1.0800 0.1830 ;
         RECT 0.9575 0.2010 0.9795 0.2870 ;
         RECT 0.9575 0.2870 0.9795 0.3010 ;
        RECT 0.9780 0.2870 1.1250 0.3010 ;
         RECT 1.1230 0.0480 1.1450 0.2010 ;
         RECT 1.1230 0.2010 1.1450 0.2870 ;
         RECT 1.1230 0.2870 1.1450 0.3010 ;
  END
END SDFFSNQ_X1

MACRO TBUF_X1
  CLASS core ;
  FOREIGN TBUF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.4620 BY 0.3840 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.1920 0.0950 0.2460 ;
         RECT 0.0730 0.2460 0.0950 0.2600 ;
        RECT 0.0930 0.2460 0.1350 0.2600 ;
        RECT 0.1350 0.2460 0.1590 0.2600 ;
         RECT 0.1570 0.1530 0.1790 0.1920 ;
         RECT 0.1570 0.1920 0.1790 0.2460 ;
         RECT 0.1570 0.2460 0.1790 0.2600 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.2830 0.1850 0.3050 0.2880 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.4085 0.0320 0.4305 0.3520 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.3860 0.3980 ;
        RECT 0.3860 0.3700 0.4690 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.4690 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0310 0.0360 0.0530 0.1560 ;
         RECT 0.0310 0.1560 0.0530 0.1700 ;
         RECT 0.0310 0.1700 0.0530 0.2090 ;
         RECT 0.0310 0.2090 0.0530 0.3430 ;
        RECT 0.0510 0.1560 0.1170 0.1700 ;
         RECT 0.1150 0.1560 0.1370 0.1700 ;
         RECT 0.1150 0.1700 0.1370 0.2090 ;
        RECT 0.0960 0.2870 0.1330 0.3010 ;
         RECT 0.1310 0.0510 0.1530 0.0650 ;
         RECT 0.1310 0.0650 0.1530 0.1150 ;
         RECT 0.1310 0.1150 0.1530 0.1290 ;
         RECT 0.1310 0.2870 0.1530 0.3010 ;
        RECT 0.1510 0.0510 0.2010 0.0650 ;
        RECT 0.1510 0.1150 0.2010 0.1290 ;
        RECT 0.1510 0.2870 0.2010 0.3010 ;
         RECT 0.1990 0.0510 0.2210 0.0650 ;
         RECT 0.1990 0.1150 0.2210 0.1290 ;
         RECT 0.1990 0.1290 0.2210 0.1570 ;
         RECT 0.1990 0.1570 0.2210 0.2870 ;
         RECT 0.1990 0.2870 0.2210 0.3010 ;
        RECT 0.2190 0.0510 0.3350 0.0650 ;
         RECT 0.3345 0.0510 0.3565 0.0650 ;
         RECT 0.3345 0.0650 0.3565 0.1150 ;
         RECT 0.3345 0.1150 0.3565 0.1290 ;
         RECT 0.3345 0.1290 0.3565 0.1570 ;
        RECT 0.0960 0.3190 0.1800 0.3330 ;
        RECT 0.1800 0.0830 0.2430 0.0970 ;
        RECT 0.1800 0.3190 0.2430 0.3330 ;
         RECT 0.2410 0.0830 0.2630 0.0970 ;
         RECT 0.2410 0.0970 0.2630 0.1880 ;
         RECT 0.2410 0.1880 0.2630 0.3190 ;
         RECT 0.2410 0.3190 0.2630 0.3330 ;
        RECT 0.2610 0.3190 0.3680 0.3330 ;
         RECT 0.3660 0.1880 0.3880 0.3190 ;
         RECT 0.3660 0.3190 0.3880 0.3330 ;
      LAYER M1 ;
         RECT 0.0310 0.0360 0.0530 0.1560 ;
         RECT 0.0310 0.1560 0.0530 0.1700 ;
         RECT 0.0310 0.1700 0.0530 0.2090 ;
         RECT 0.0310 0.2090 0.0530 0.3430 ;
        RECT 0.0510 0.1560 0.1170 0.1700 ;
         RECT 0.1150 0.1560 0.1370 0.1700 ;
         RECT 0.1150 0.1700 0.1370 0.2090 ;
        RECT 0.0960 0.2870 0.1330 0.3010 ;
         RECT 0.1310 0.0510 0.1530 0.0650 ;
         RECT 0.1310 0.0650 0.1530 0.1150 ;
         RECT 0.1310 0.1150 0.1530 0.1290 ;
         RECT 0.1310 0.2870 0.1530 0.3010 ;
        RECT 0.1510 0.0510 0.2010 0.0650 ;
        RECT 0.1510 0.1150 0.2010 0.1290 ;
        RECT 0.1510 0.2870 0.2010 0.3010 ;
         RECT 0.1990 0.0510 0.2210 0.0650 ;
         RECT 0.1990 0.1150 0.2210 0.1290 ;
         RECT 0.1990 0.1290 0.2210 0.1570 ;
         RECT 0.1990 0.1570 0.2210 0.2870 ;
         RECT 0.1990 0.2870 0.2210 0.3010 ;
        RECT 0.2190 0.0510 0.3350 0.0650 ;
         RECT 0.3345 0.0510 0.3565 0.0650 ;
         RECT 0.3345 0.0650 0.3565 0.1150 ;
         RECT 0.3345 0.1150 0.3565 0.1290 ;
         RECT 0.3345 0.1290 0.3565 0.1570 ;
        RECT 0.0960 0.3190 0.1800 0.3330 ;
        RECT 0.1800 0.0830 0.2430 0.0970 ;
        RECT 0.1800 0.3190 0.2430 0.3330 ;
         RECT 0.2410 0.0830 0.2630 0.0970 ;
         RECT 0.2410 0.0970 0.2630 0.1880 ;
         RECT 0.2410 0.1880 0.2630 0.3190 ;
         RECT 0.2410 0.3190 0.2630 0.3330 ;
        RECT 0.2610 0.3190 0.3680 0.3330 ;
         RECT 0.3660 0.1880 0.3880 0.3190 ;
         RECT 0.3660 0.3190 0.3880 0.3330 ;
  END
END TBUF_X1

MACRO TBUF_X2
  CLASS core ;
  FOREIGN TBUF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.5040 BY 0.3840 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.1920 0.0950 0.2520 ;
         RECT 0.0730 0.2520 0.0950 0.2660 ;
        RECT 0.0930 0.2520 0.1350 0.2660 ;
        RECT 0.1350 0.2520 0.1590 0.2660 ;
         RECT 0.1570 0.1530 0.1790 0.1920 ;
         RECT 0.1570 0.1920 0.1790 0.2520 ;
         RECT 0.1570 0.2520 0.1790 0.2660 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.2830 0.1910 0.3050 0.2880 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.4085 0.0350 0.4305 0.3480 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.3480 0.3980 ;
        RECT 0.3480 0.3700 0.5110 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.5110 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0310 0.0360 0.0530 0.1560 ;
         RECT 0.0310 0.1560 0.0530 0.1700 ;
         RECT 0.0310 0.1700 0.0530 0.2020 ;
         RECT 0.0310 0.2020 0.0530 0.3060 ;
        RECT 0.0510 0.1560 0.1170 0.1700 ;
         RECT 0.1150 0.1560 0.1370 0.1700 ;
         RECT 0.1150 0.1700 0.1370 0.2020 ;
        RECT 0.0960 0.2840 0.1330 0.3010 ;
         RECT 0.1310 0.0510 0.1530 0.0650 ;
         RECT 0.1310 0.0650 0.1530 0.1150 ;
         RECT 0.1310 0.1150 0.1530 0.1290 ;
         RECT 0.1310 0.2840 0.1530 0.3010 ;
        RECT 0.1510 0.0510 0.2010 0.0650 ;
        RECT 0.1510 0.1150 0.2010 0.1290 ;
        RECT 0.1510 0.2840 0.2010 0.3010 ;
         RECT 0.1990 0.0510 0.2210 0.0650 ;
         RECT 0.1990 0.1150 0.2210 0.1290 ;
         RECT 0.1990 0.1290 0.2210 0.1570 ;
         RECT 0.1990 0.1570 0.2210 0.2840 ;
         RECT 0.1990 0.2840 0.2210 0.3010 ;
        RECT 0.2190 0.0510 0.3160 0.0650 ;
         RECT 0.3155 0.0510 0.3375 0.0650 ;
         RECT 0.3155 0.0650 0.3375 0.1150 ;
         RECT 0.3155 0.1150 0.3375 0.1290 ;
         RECT 0.3155 0.1290 0.3375 0.1570 ;
        RECT 0.0960 0.3190 0.1800 0.3330 ;
        RECT 0.1800 0.0830 0.2430 0.0970 ;
        RECT 0.1800 0.3190 0.2430 0.3330 ;
         RECT 0.2410 0.0830 0.2630 0.0970 ;
         RECT 0.2410 0.0970 0.2630 0.2220 ;
         RECT 0.2410 0.2220 0.2630 0.3190 ;
         RECT 0.2410 0.3190 0.2630 0.3330 ;
        RECT 0.2610 0.3190 0.3270 0.3330 ;
         RECT 0.3265 0.2220 0.3485 0.3190 ;
         RECT 0.3265 0.3190 0.3485 0.3330 ;
      LAYER M1 ;
         RECT 0.0310 0.0360 0.0530 0.1560 ;
         RECT 0.0310 0.1560 0.0530 0.1700 ;
         RECT 0.0310 0.1700 0.0530 0.2020 ;
         RECT 0.0310 0.2020 0.0530 0.3060 ;
        RECT 0.0510 0.1560 0.1170 0.1700 ;
         RECT 0.1150 0.1560 0.1370 0.1700 ;
         RECT 0.1150 0.1700 0.1370 0.2020 ;
        RECT 0.0960 0.2840 0.1330 0.3010 ;
         RECT 0.1310 0.0510 0.1530 0.0650 ;
         RECT 0.1310 0.0650 0.1530 0.1150 ;
         RECT 0.1310 0.1150 0.1530 0.1290 ;
         RECT 0.1310 0.2840 0.1530 0.3010 ;
        RECT 0.1510 0.0510 0.2010 0.0650 ;
        RECT 0.1510 0.1150 0.2010 0.1290 ;
        RECT 0.1510 0.2840 0.2010 0.3010 ;
         RECT 0.1990 0.0510 0.2210 0.0650 ;
         RECT 0.1990 0.1150 0.2210 0.1290 ;
         RECT 0.1990 0.1290 0.2210 0.1570 ;
         RECT 0.1990 0.1570 0.2210 0.2840 ;
         RECT 0.1990 0.2840 0.2210 0.3010 ;
        RECT 0.2190 0.0510 0.3160 0.0650 ;
         RECT 0.3155 0.0510 0.3375 0.0650 ;
         RECT 0.3155 0.0650 0.3375 0.1150 ;
         RECT 0.3155 0.1150 0.3375 0.1290 ;
         RECT 0.3155 0.1290 0.3375 0.1570 ;
        RECT 0.0960 0.3190 0.1800 0.3330 ;
        RECT 0.1800 0.0830 0.2430 0.0970 ;
        RECT 0.1800 0.3190 0.2430 0.3330 ;
         RECT 0.2410 0.0830 0.2630 0.0970 ;
         RECT 0.2410 0.0970 0.2630 0.2220 ;
         RECT 0.2410 0.2220 0.2630 0.3190 ;
         RECT 0.2410 0.3190 0.2630 0.3330 ;
        RECT 0.2610 0.3190 0.3270 0.3330 ;
         RECT 0.3265 0.2220 0.3485 0.3190 ;
         RECT 0.3265 0.3190 0.3485 0.3330 ;
  END
END TBUF_X2

MACRO TBUF_X4
  CLASS core ;
  FOREIGN TBUF_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.6300 BY 0.3840 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.1920 0.0950 0.2420 ;
         RECT 0.0730 0.2420 0.0950 0.2560 ;
        RECT 0.0930 0.2420 0.1350 0.2560 ;
        RECT 0.1350 0.2420 0.1590 0.2560 ;
         RECT 0.1570 0.1530 0.1790 0.1920 ;
         RECT 0.1570 0.1920 0.1790 0.2420 ;
         RECT 0.1570 0.2420 0.1790 0.2560 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.2830 0.1730 0.3050 0.2970 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.4505 0.0320 0.4725 0.1120 ;
         RECT 0.4505 0.1120 0.4725 0.1280 ;
         RECT 0.4505 0.2560 0.4725 0.2700 ;
         RECT 0.4505 0.2700 0.4725 0.2850 ;
         RECT 0.4505 0.2850 0.4725 0.3520 ;
        RECT 0.4720 0.1120 0.5330 0.1280 ;
        RECT 0.4720 0.2560 0.5330 0.2700 ;
         RECT 0.5225 0.0320 0.5445 0.1120 ;
         RECT 0.5225 0.1120 0.5445 0.1280 ;
         RECT 0.5225 0.2560 0.5445 0.2700 ;
         RECT 0.5235 0.0320 0.5455 0.1120 ;
         RECT 0.5235 0.1120 0.5455 0.1280 ;
         RECT 0.5235 0.2560 0.5455 0.2700 ;
         RECT 0.5315 0.0320 0.5535 0.1120 ;
         RECT 0.5315 0.1120 0.5535 0.1280 ;
         RECT 0.5315 0.2560 0.5535 0.2700 ;
         RECT 0.5315 0.2700 0.5535 0.2850 ;
         RECT 0.5315 0.2850 0.5535 0.3520 ;
         RECT 0.5420 0.0320 0.5640 0.1120 ;
         RECT 0.5420 0.1120 0.5640 0.1280 ;
         RECT 0.5420 0.2560 0.5640 0.2700 ;
         RECT 0.5420 0.2700 0.5640 0.2850 ;
         RECT 0.5420 0.2850 0.5640 0.3520 ;
         RECT 0.5460 0.0320 0.5680 0.1120 ;
         RECT 0.5460 0.1120 0.5680 0.1280 ;
         RECT 0.5460 0.2560 0.5680 0.2700 ;
         RECT 0.5460 0.2700 0.5680 0.2850 ;
         RECT 0.5575 0.1120 0.5795 0.1280 ;
         RECT 0.5575 0.2560 0.5795 0.2700 ;
         RECT 0.5575 0.2700 0.5795 0.2850 ;
         RECT 0.5770 0.1120 0.5990 0.1280 ;
         RECT 0.5770 0.1280 0.5990 0.2560 ;
         RECT 0.5770 0.2560 0.5990 0.2700 ;
         RECT 0.5770 0.2700 0.5990 0.2850 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.5340 0.3980 ;
         RECT 0.5310 0.3700 0.5530 0.3980 ;
        RECT 0.5500 0.3700 0.6370 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.6370 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.0540 0.3190 0.1800 0.3330 ;
        RECT 0.1800 0.0830 0.2430 0.0970 ;
        RECT 0.1800 0.3190 0.2430 0.3330 ;
         RECT 0.2410 0.0830 0.2630 0.0970 ;
         RECT 0.2410 0.0970 0.2630 0.1940 ;
         RECT 0.2410 0.1940 0.2630 0.2070 ;
         RECT 0.2410 0.2070 0.2630 0.2290 ;
         RECT 0.2410 0.2290 0.2630 0.3190 ;
         RECT 0.2410 0.3190 0.2630 0.3330 ;
        RECT 0.2610 0.3190 0.3450 0.3330 ;
        RECT 0.3450 0.1940 0.3820 0.2070 ;
        RECT 0.3450 0.2070 0.3820 0.2290 ;
        RECT 0.3450 0.2290 0.3820 0.3190 ;
        RECT 0.3450 0.3190 0.3820 0.3330 ;
        RECT 0.3820 0.2070 0.5340 0.2290 ;
         RECT 0.0310 0.0480 0.0530 0.1560 ;
         RECT 0.0310 0.1560 0.0530 0.1700 ;
         RECT 0.0310 0.1700 0.0530 0.2020 ;
         RECT 0.0310 0.2020 0.0530 0.2970 ;
        RECT 0.0510 0.1560 0.1170 0.1700 ;
         RECT 0.1150 0.1560 0.1370 0.1700 ;
         RECT 0.1150 0.1700 0.1370 0.2020 ;
        RECT 0.0960 0.2840 0.1330 0.3010 ;
         RECT 0.1310 0.0510 0.1530 0.0650 ;
         RECT 0.1310 0.0650 0.1530 0.1150 ;
         RECT 0.1310 0.1150 0.1530 0.1290 ;
         RECT 0.1310 0.2840 0.1530 0.3010 ;
        RECT 0.1510 0.0510 0.2010 0.0650 ;
        RECT 0.1510 0.1150 0.2010 0.1290 ;
        RECT 0.1510 0.2840 0.2010 0.3010 ;
         RECT 0.1990 0.0510 0.2210 0.0650 ;
         RECT 0.1990 0.1150 0.2210 0.1290 ;
         RECT 0.1990 0.1290 0.2210 0.1460 ;
         RECT 0.1990 0.1460 0.2210 0.1600 ;
         RECT 0.1990 0.1600 0.2210 0.1760 ;
         RECT 0.1990 0.1760 0.2210 0.2840 ;
         RECT 0.1990 0.2840 0.2210 0.3010 ;
        RECT 0.2190 0.0510 0.3450 0.0650 ;
        RECT 0.3450 0.0510 0.3820 0.0650 ;
        RECT 0.3450 0.0650 0.3820 0.1150 ;
        RECT 0.3450 0.1150 0.3820 0.1290 ;
        RECT 0.3450 0.1290 0.3820 0.1460 ;
        RECT 0.3450 0.1460 0.3820 0.1600 ;
        RECT 0.3450 0.1600 0.3820 0.1760 ;
        RECT 0.3820 0.1460 0.5500 0.1600 ;
      LAYER M1 ;
        RECT 0.0540 0.3190 0.1800 0.3330 ;
        RECT 0.1800 0.0830 0.2430 0.0970 ;
        RECT 0.1800 0.3190 0.2430 0.3330 ;
         RECT 0.2410 0.0830 0.2630 0.0970 ;
         RECT 0.2410 0.0970 0.2630 0.1940 ;
         RECT 0.2410 0.1940 0.2630 0.2070 ;
         RECT 0.2410 0.2070 0.2630 0.2290 ;
         RECT 0.2410 0.2290 0.2630 0.3190 ;
         RECT 0.2410 0.3190 0.2630 0.3330 ;
        RECT 0.2610 0.3190 0.3450 0.3330 ;
        RECT 0.3450 0.1940 0.3820 0.2070 ;
        RECT 0.3450 0.2070 0.3820 0.2290 ;
        RECT 0.3450 0.2290 0.3820 0.3190 ;
        RECT 0.3450 0.3190 0.3820 0.3330 ;
        RECT 0.3820 0.2070 0.5340 0.2290 ;
         RECT 0.0310 0.0480 0.0530 0.1560 ;
         RECT 0.0310 0.1560 0.0530 0.1700 ;
         RECT 0.0310 0.1700 0.0530 0.2020 ;
         RECT 0.0310 0.2020 0.0530 0.2970 ;
        RECT 0.0510 0.1560 0.1170 0.1700 ;
         RECT 0.1150 0.1560 0.1370 0.1700 ;
         RECT 0.1150 0.1700 0.1370 0.2020 ;
        RECT 0.0960 0.2840 0.1330 0.3010 ;
         RECT 0.1310 0.0510 0.1530 0.0650 ;
         RECT 0.1310 0.0650 0.1530 0.1150 ;
         RECT 0.1310 0.1150 0.1530 0.1290 ;
         RECT 0.1310 0.2840 0.1530 0.3010 ;
        RECT 0.1510 0.0510 0.2010 0.0650 ;
        RECT 0.1510 0.1150 0.2010 0.1290 ;
        RECT 0.1510 0.2840 0.2010 0.3010 ;
         RECT 0.1990 0.0510 0.2210 0.0650 ;
         RECT 0.1990 0.1150 0.2210 0.1290 ;
         RECT 0.1990 0.1290 0.2210 0.1460 ;
         RECT 0.1990 0.1460 0.2210 0.1600 ;
         RECT 0.1990 0.1600 0.2210 0.1760 ;
         RECT 0.1990 0.1760 0.2210 0.2840 ;
         RECT 0.1990 0.2840 0.2210 0.3010 ;
        RECT 0.2190 0.0510 0.3450 0.0650 ;
        RECT 0.3450 0.0510 0.3820 0.0650 ;
        RECT 0.3450 0.0650 0.3820 0.1150 ;
        RECT 0.3450 0.1150 0.3820 0.1290 ;
        RECT 0.3450 0.1290 0.3820 0.1460 ;
        RECT 0.3450 0.1460 0.3820 0.1600 ;
        RECT 0.3450 0.1600 0.3820 0.1760 ;
        RECT 0.3820 0.1460 0.5500 0.1600 ;
  END
END TBUF_X4

MACRO TBUF_X8
  CLASS core ;
  FOREIGN TBUF_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.8820 BY 0.3840 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.1920 0.0950 0.2420 ;
         RECT 0.0730 0.2420 0.0950 0.2560 ;
        RECT 0.0930 0.2420 0.1460 0.2560 ;
        RECT 0.1460 0.2420 0.2010 0.2560 ;
         RECT 0.1990 0.1600 0.2210 0.1920 ;
         RECT 0.1990 0.1920 0.2210 0.2420 ;
         RECT 0.1990 0.2420 0.2210 0.2560 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.3250 0.1730 0.3470 0.2010 ;
         RECT 0.3250 0.2010 0.3470 0.2170 ;
         RECT 0.3250 0.2170 0.3470 0.2880 ;
        RECT 0.3450 0.2010 0.4080 0.2170 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.5345 0.0320 0.5565 0.0660 ;
         RECT 0.5345 0.0660 0.5565 0.0800 ;
         RECT 0.5345 0.0800 0.5565 0.0960 ;
         RECT 0.5345 0.2600 0.5565 0.2880 ;
         RECT 0.5345 0.2880 0.5565 0.2890 ;
         RECT 0.5345 0.2890 0.5565 0.3520 ;
        RECT 0.5560 0.0800 0.7760 0.0960 ;
        RECT 0.5560 0.2600 0.7760 0.2880 ;
         RECT 0.7700 0.0800 0.7920 0.0960 ;
         RECT 0.7700 0.2600 0.7920 0.2880 ;
         RECT 0.7760 0.0800 0.7980 0.0960 ;
         RECT 0.7760 0.2600 0.7980 0.2880 ;
         RECT 0.7870 0.0320 0.8090 0.0660 ;
         RECT 0.7870 0.0660 0.8090 0.0800 ;
         RECT 0.7870 0.0800 0.8090 0.0960 ;
         RECT 0.7870 0.2600 0.8090 0.2880 ;
         RECT 0.7870 0.2880 0.8090 0.2890 ;
         RECT 0.7870 0.2890 0.8090 0.3520 ;
        RECT 0.8080 0.0660 0.8310 0.0800 ;
        RECT 0.8080 0.0800 0.8310 0.0960 ;
        RECT 0.8080 0.2600 0.8310 0.2880 ;
        RECT 0.8080 0.2880 0.8310 0.2890 ;
         RECT 0.8290 0.0660 0.8510 0.0800 ;
         RECT 0.8290 0.0800 0.8510 0.0960 ;
         RECT 0.8290 0.0960 0.8510 0.2600 ;
         RECT 0.8290 0.2600 0.8510 0.2880 ;
         RECT 0.8290 0.2880 0.8510 0.2890 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.7760 0.3980 ;
         RECT 0.7700 0.3700 0.7920 0.3980 ;
        RECT 0.7860 0.3700 0.8890 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.8890 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0310 0.0360 0.0530 0.1560 ;
         RECT 0.0310 0.1560 0.0530 0.1700 ;
         RECT 0.0310 0.1700 0.0530 0.2150 ;
         RECT 0.0310 0.2150 0.0530 0.3190 ;
        RECT 0.0510 0.1560 0.1170 0.1700 ;
        RECT 0.1170 0.1560 0.1460 0.1700 ;
        RECT 0.1170 0.1700 0.1460 0.2150 ;
        RECT 0.0960 0.2870 0.1330 0.3010 ;
         RECT 0.1310 0.0510 0.1530 0.0650 ;
         RECT 0.1310 0.0650 0.1530 0.1150 ;
         RECT 0.1310 0.1150 0.1530 0.1290 ;
         RECT 0.1310 0.2870 0.1530 0.3010 ;
        RECT 0.1510 0.0510 0.2430 0.0650 ;
        RECT 0.1510 0.1150 0.2430 0.1290 ;
        RECT 0.1510 0.2870 0.2430 0.3010 ;
         RECT 0.2410 0.0510 0.2630 0.0650 ;
         RECT 0.2410 0.1150 0.2630 0.1290 ;
         RECT 0.2410 0.1290 0.2630 0.1430 ;
         RECT 0.2410 0.1430 0.2630 0.1710 ;
         RECT 0.2410 0.1710 0.2630 0.2870 ;
         RECT 0.2410 0.2870 0.2630 0.3010 ;
        RECT 0.2610 0.0510 0.4530 0.0650 ;
         RECT 0.4510 0.0510 0.4730 0.0650 ;
         RECT 0.4510 0.0650 0.4730 0.1150 ;
         RECT 0.4510 0.1150 0.4730 0.1290 ;
         RECT 0.4510 0.1290 0.4730 0.1430 ;
         RECT 0.4510 0.1430 0.4730 0.1710 ;
        RECT 0.4710 0.1290 0.7860 0.1430 ;
        RECT 0.0800 0.3190 0.1800 0.3330 ;
        RECT 0.1800 0.0830 0.2850 0.0970 ;
        RECT 0.1800 0.3190 0.2850 0.3330 ;
         RECT 0.2830 0.0830 0.3050 0.0970 ;
         RECT 0.2830 0.0970 0.3050 0.1930 ;
         RECT 0.2830 0.1930 0.3050 0.2020 ;
         RECT 0.2830 0.2020 0.3050 0.2300 ;
         RECT 0.2830 0.2300 0.3050 0.3190 ;
         RECT 0.2830 0.3190 0.3050 0.3330 ;
        RECT 0.3030 0.3190 0.4330 0.3330 ;
        RECT 0.4330 0.1930 0.4710 0.2020 ;
        RECT 0.4330 0.2020 0.4710 0.2300 ;
        RECT 0.4330 0.2300 0.4710 0.3190 ;
        RECT 0.4330 0.3190 0.4710 0.3330 ;
        RECT 0.4710 0.2020 0.7760 0.2300 ;
      LAYER M1 ;
         RECT 0.0310 0.0360 0.0530 0.1560 ;
         RECT 0.0310 0.1560 0.0530 0.1700 ;
         RECT 0.0310 0.1700 0.0530 0.2150 ;
         RECT 0.0310 0.2150 0.0530 0.3190 ;
        RECT 0.0510 0.1560 0.1170 0.1700 ;
        RECT 0.1170 0.1560 0.1460 0.1700 ;
        RECT 0.1170 0.1700 0.1460 0.2150 ;
        RECT 0.0960 0.2870 0.1330 0.3010 ;
         RECT 0.1310 0.0510 0.1530 0.0650 ;
         RECT 0.1310 0.0650 0.1530 0.1150 ;
         RECT 0.1310 0.1150 0.1530 0.1290 ;
         RECT 0.1310 0.2870 0.1530 0.3010 ;
        RECT 0.1510 0.0510 0.2430 0.0650 ;
        RECT 0.1510 0.1150 0.2430 0.1290 ;
        RECT 0.1510 0.2870 0.2430 0.3010 ;
         RECT 0.2410 0.0510 0.2630 0.0650 ;
         RECT 0.2410 0.1150 0.2630 0.1290 ;
         RECT 0.2410 0.1290 0.2630 0.1430 ;
         RECT 0.2410 0.1430 0.2630 0.1710 ;
         RECT 0.2410 0.1710 0.2630 0.2870 ;
         RECT 0.2410 0.2870 0.2630 0.3010 ;
        RECT 0.2610 0.0510 0.4530 0.0650 ;
         RECT 0.4510 0.0510 0.4730 0.0650 ;
         RECT 0.4510 0.0650 0.4730 0.1150 ;
         RECT 0.4510 0.1150 0.4730 0.1290 ;
         RECT 0.4510 0.1290 0.4730 0.1430 ;
         RECT 0.4510 0.1430 0.4730 0.1710 ;
        RECT 0.4710 0.1290 0.7860 0.1430 ;
        RECT 0.0800 0.3190 0.1800 0.3330 ;
        RECT 0.1800 0.0830 0.2850 0.0970 ;
        RECT 0.1800 0.3190 0.2850 0.3330 ;
         RECT 0.2830 0.0830 0.3050 0.0970 ;
         RECT 0.2830 0.0970 0.3050 0.1930 ;
         RECT 0.2830 0.1930 0.3050 0.2020 ;
         RECT 0.2830 0.2020 0.3050 0.2300 ;
         RECT 0.2830 0.2300 0.3050 0.3190 ;
         RECT 0.2830 0.3190 0.3050 0.3330 ;
        RECT 0.3030 0.3190 0.4330 0.3330 ;
        RECT 0.4330 0.1930 0.4710 0.2020 ;
        RECT 0.4330 0.2020 0.4710 0.2300 ;
        RECT 0.4330 0.2300 0.4710 0.3190 ;
        RECT 0.4330 0.3190 0.4710 0.3330 ;
        RECT 0.4710 0.2020 0.7760 0.2300 ;
  END
END TBUF_X8

MACRO TBUF_X12
  CLASS core ;
  FOREIGN TBUF_X12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 1.1340 BY 0.3840 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.1920 0.0950 0.2550 ;
         RECT 0.0730 0.2550 0.0950 0.2690 ;
        RECT 0.0930 0.2550 0.1350 0.2690 ;
        RECT 0.1350 0.2550 0.1590 0.2690 ;
         RECT 0.1570 0.1530 0.1790 0.1920 ;
         RECT 0.1570 0.1920 0.1790 0.2550 ;
         RECT 0.1570 0.2550 0.1790 0.2690 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.2850 0.2010 0.3270 0.2240 ;
         RECT 0.3250 0.1730 0.3470 0.2010 ;
         RECT 0.3250 0.2010 0.3470 0.2240 ;
        RECT 0.3450 0.2010 0.4110 0.2240 ;
         RECT 0.4090 0.2010 0.4310 0.2240 ;
         RECT 0.4090 0.2240 0.4310 0.2880 ;
        RECT 0.4290 0.2010 0.4660 0.2240 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 1.1050 0.3980 ;
        RECT 1.1050 0.3700 1.1410 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 1.1410 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.0960 0.3190 0.1800 0.3330 ;
        RECT 0.1800 0.0830 0.2430 0.0970 ;
        RECT 0.1800 0.3190 0.2430 0.3330 ;
         RECT 0.2410 0.0830 0.2630 0.0970 ;
         RECT 0.2410 0.0970 0.2630 0.1780 ;
         RECT 0.2410 0.1780 0.2630 0.1890 ;
         RECT 0.2410 0.1890 0.2630 0.2130 ;
         RECT 0.2410 0.2130 0.2630 0.3190 ;
         RECT 0.2410 0.3190 0.2630 0.3330 ;
        RECT 0.2610 0.3190 0.5140 0.3330 ;
        RECT 0.5140 0.1780 0.5510 0.1890 ;
        RECT 0.5140 0.1890 0.5510 0.2130 ;
        RECT 0.5140 0.2130 0.5510 0.3190 ;
        RECT 0.5140 0.3190 0.5510 0.3330 ;
        RECT 0.5510 0.1890 1.0220 0.2130 ;
        RECT 0.5790 0.0510 0.6110 0.0650 ;
        RECT 0.6110 0.0510 0.6490 0.0650 ;
        RECT 0.6110 0.2660 0.6490 0.2820 ;
        RECT 0.6110 0.2820 0.6490 0.3100 ;
        RECT 0.6490 0.0510 1.0320 0.0650 ;
        RECT 0.6490 0.2660 1.0320 0.2820 ;
         RECT 1.0255 0.0360 1.0475 0.0510 ;
         RECT 1.0255 0.0510 1.0475 0.0650 ;
         RECT 1.0255 0.2660 1.0475 0.2820 ;
         RECT 1.0390 0.0360 1.0610 0.0510 ;
         RECT 1.0390 0.0510 1.0610 0.0650 ;
         RECT 1.0390 0.2660 1.0610 0.2820 ;
         RECT 1.0390 0.2820 1.0610 0.3100 ;
         RECT 1.0390 0.3100 1.0610 0.3120 ;
         RECT 1.0525 0.0360 1.0745 0.0510 ;
         RECT 1.0525 0.0510 1.0745 0.0650 ;
         RECT 1.0525 0.2660 1.0745 0.2820 ;
         RECT 1.0575 0.0510 1.0795 0.0650 ;
         RECT 1.0575 0.2660 1.0795 0.2820 ;
        RECT 1.0690 0.0510 1.1050 0.0650 ;
        RECT 1.0690 0.0650 1.1050 0.2660 ;
        RECT 1.0690 0.2660 1.1050 0.2820 ;
         RECT 0.0310 0.0870 0.0530 0.1560 ;
         RECT 0.0310 0.1560 0.0530 0.1700 ;
         RECT 0.0310 0.1700 0.0530 0.2020 ;
         RECT 0.0310 0.2020 0.0530 0.3360 ;
        RECT 0.0510 0.1560 0.1170 0.1700 ;
         RECT 0.1150 0.1560 0.1370 0.1700 ;
         RECT 0.1150 0.1700 0.1370 0.2020 ;
         RECT 0.0835 0.0510 0.1055 0.0650 ;
         RECT 0.0835 0.0650 0.1055 0.1150 ;
         RECT 0.0835 0.1150 0.1055 0.1250 ;
         RECT 0.0835 0.1250 0.1055 0.1290 ;
         RECT 0.0930 0.0510 0.1150 0.0650 ;
         RECT 0.0930 0.0650 0.1150 0.1150 ;
         RECT 0.0930 0.1150 0.1150 0.1250 ;
         RECT 0.0930 0.1250 0.1150 0.1290 ;
         RECT 0.0930 0.2870 0.1150 0.3010 ;
        RECT 0.1120 0.0510 0.2010 0.0650 ;
        RECT 0.1120 0.1150 0.2010 0.1250 ;
        RECT 0.1120 0.1250 0.2010 0.1290 ;
        RECT 0.1120 0.2870 0.2010 0.3010 ;
         RECT 0.1990 0.0510 0.2210 0.0650 ;
         RECT 0.1990 0.1150 0.2210 0.1250 ;
         RECT 0.1990 0.1250 0.2210 0.1290 ;
         RECT 0.1990 0.1290 0.2210 0.1470 ;
         RECT 0.1990 0.1470 0.2210 0.2870 ;
         RECT 0.1990 0.2870 0.2210 0.3010 ;
        RECT 0.2190 0.0510 0.5130 0.0650 ;
         RECT 0.5125 0.0510 0.5345 0.0650 ;
         RECT 0.5125 0.0650 0.5345 0.1150 ;
         RECT 0.5125 0.1150 0.5345 0.1250 ;
         RECT 0.5125 0.1250 0.5345 0.1290 ;
         RECT 0.5125 0.1290 0.5345 0.1470 ;
        RECT 0.5340 0.1250 1.0450 0.1290 ;
        RECT 0.5340 0.1290 1.0450 0.1470 ;
      LAYER M1 ;
        RECT 0.0960 0.3190 0.1800 0.3330 ;
        RECT 0.1800 0.0830 0.2430 0.0970 ;
        RECT 0.1800 0.3190 0.2430 0.3330 ;
         RECT 0.2410 0.0830 0.2630 0.0970 ;
         RECT 0.2410 0.0970 0.2630 0.1780 ;
         RECT 0.2410 0.1780 0.2630 0.1890 ;
         RECT 0.2410 0.1890 0.2630 0.2130 ;
         RECT 0.2410 0.2130 0.2630 0.3190 ;
         RECT 0.2410 0.3190 0.2630 0.3330 ;
        RECT 0.2610 0.3190 0.5140 0.3330 ;
        RECT 0.5140 0.1780 0.5510 0.1890 ;
        RECT 0.5140 0.1890 0.5510 0.2130 ;
        RECT 0.5140 0.2130 0.5510 0.3190 ;
        RECT 0.5140 0.3190 0.5510 0.3330 ;
        RECT 0.5510 0.1890 1.0220 0.2130 ;
        RECT 0.5790 0.0510 0.6110 0.0650 ;
        RECT 0.6110 0.0510 0.6490 0.0650 ;
        RECT 0.6110 0.2660 0.6490 0.2820 ;
        RECT 0.6110 0.2820 0.6490 0.3100 ;
        RECT 0.6490 0.0510 1.0320 0.0650 ;
        RECT 0.6490 0.2660 1.0320 0.2820 ;
         RECT 1.0255 0.0360 1.0475 0.0510 ;
         RECT 1.0255 0.0510 1.0475 0.0650 ;
         RECT 1.0255 0.2660 1.0475 0.2820 ;
         RECT 1.0390 0.0360 1.0610 0.0510 ;
         RECT 1.0390 0.0510 1.0610 0.0650 ;
         RECT 1.0390 0.2660 1.0610 0.2820 ;
         RECT 1.0390 0.2820 1.0610 0.3100 ;
         RECT 1.0390 0.3100 1.0610 0.3120 ;
         RECT 1.0525 0.0360 1.0745 0.0510 ;
         RECT 1.0525 0.0510 1.0745 0.0650 ;
         RECT 1.0525 0.2660 1.0745 0.2820 ;
         RECT 1.0575 0.0510 1.0795 0.0650 ;
         RECT 1.0575 0.2660 1.0795 0.2820 ;
        RECT 1.0690 0.0510 1.1050 0.0650 ;
        RECT 1.0690 0.0650 1.1050 0.2660 ;
        RECT 1.0690 0.2660 1.1050 0.2820 ;
         RECT 0.0310 0.0870 0.0530 0.1560 ;
         RECT 0.0310 0.1560 0.0530 0.1700 ;
         RECT 0.0310 0.1700 0.0530 0.2020 ;
         RECT 0.0310 0.2020 0.0530 0.3360 ;
        RECT 0.0510 0.1560 0.1170 0.1700 ;
         RECT 0.1150 0.1560 0.1370 0.1700 ;
         RECT 0.1150 0.1700 0.1370 0.2020 ;
         RECT 0.0835 0.0510 0.1055 0.0650 ;
         RECT 0.0835 0.0650 0.1055 0.1150 ;
         RECT 0.0835 0.1150 0.1055 0.1250 ;
         RECT 0.0835 0.1250 0.1055 0.1290 ;
         RECT 0.0930 0.0510 0.1150 0.0650 ;
         RECT 0.0930 0.0650 0.1150 0.1150 ;
         RECT 0.0930 0.1150 0.1150 0.1250 ;
         RECT 0.0930 0.1250 0.1150 0.1290 ;
         RECT 0.0930 0.2870 0.1150 0.3010 ;
        RECT 0.1120 0.0510 0.2010 0.0650 ;
        RECT 0.1120 0.1150 0.2010 0.1250 ;
        RECT 0.1120 0.1250 0.2010 0.1290 ;
        RECT 0.1120 0.2870 0.2010 0.3010 ;
         RECT 0.1990 0.0510 0.2210 0.0650 ;
         RECT 0.1990 0.1150 0.2210 0.1250 ;
         RECT 0.1990 0.1250 0.2210 0.1290 ;
         RECT 0.1990 0.1290 0.2210 0.1470 ;
         RECT 0.1990 0.1470 0.2210 0.2870 ;
         RECT 0.1990 0.2870 0.2210 0.3010 ;
        RECT 0.2190 0.0510 0.5130 0.0650 ;
         RECT 0.5125 0.0510 0.5345 0.0650 ;
         RECT 0.5125 0.0650 0.5345 0.1150 ;
         RECT 0.5125 0.1150 0.5345 0.1250 ;
         RECT 0.5125 0.1250 0.5345 0.1290 ;
         RECT 0.5125 0.1290 0.5345 0.1470 ;
        RECT 0.5340 0.1250 1.0450 0.1290 ;
        RECT 0.5340 0.1290 1.0450 0.1470 ;
  END
END TBUF_X12

MACRO TBUF_X16
  CLASS core ;
  FOREIGN TBUF_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 1.3860 BY 0.3840 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0730 0.1950 0.0950 0.2430 ;
         RECT 0.0730 0.2430 0.0950 0.2570 ;
         RECT 0.0925 0.2430 0.1145 0.2570 ;
        RECT 0.1140 0.2430 0.1580 0.2570 ;
         RECT 0.1575 0.1600 0.1795 0.1950 ;
         RECT 0.1575 0.1950 0.1795 0.2430 ;
         RECT 0.1575 0.2430 0.1795 0.2570 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.3030 0.2010 0.3690 0.2240 ;
         RECT 0.3670 0.1730 0.3890 0.2010 ;
         RECT 0.3670 0.2010 0.3890 0.2240 ;
        RECT 0.3870 0.2010 0.4530 0.2240 ;
         RECT 0.4510 0.2010 0.4730 0.2240 ;
         RECT 0.4510 0.2240 0.4730 0.2880 ;
        RECT 0.4710 0.2010 0.5920 0.2240 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.7030 0.0320 0.7250 0.0710 ;
         RECT 0.7030 0.0710 0.7250 0.1000 ;
         RECT 0.7030 0.2600 0.7250 0.2880 ;
         RECT 0.7030 0.2880 0.7250 0.3520 ;
        RECT 0.7240 0.0710 1.2920 0.1000 ;
        RECT 0.7240 0.2600 1.2920 0.2880 ;
         RECT 1.2845 0.0320 1.3065 0.0710 ;
         RECT 1.2845 0.0710 1.3065 0.1000 ;
         RECT 1.2845 0.2600 1.3065 0.2880 ;
         RECT 1.2845 0.2880 1.3065 0.3520 ;
         RECT 1.2940 0.0320 1.3160 0.0710 ;
         RECT 1.2940 0.0710 1.3160 0.1000 ;
         RECT 1.2940 0.2600 1.3160 0.2880 ;
         RECT 1.2940 0.2880 1.3160 0.3520 ;
         RECT 1.3005 0.0320 1.3225 0.0710 ;
         RECT 1.3005 0.0710 1.3225 0.1000 ;
         RECT 1.3005 0.2600 1.3225 0.2880 ;
         RECT 1.3005 0.2880 1.3225 0.3520 ;
        RECT 1.3120 0.0710 1.3350 0.1000 ;
        RECT 1.3120 0.2600 1.3350 0.2880 ;
         RECT 1.3330 0.0710 1.3550 0.1000 ;
         RECT 1.3330 0.1000 1.3550 0.2600 ;
         RECT 1.3330 0.2600 1.3550 0.2880 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 1.2990 0.3980 ;
         RECT 1.2940 0.3700 1.3160 0.3980 ;
        RECT 1.3110 0.3700 1.3930 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 1.3930 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0310 0.0360 0.0530 0.1310 ;
         RECT 0.0310 0.1310 0.0530 0.1450 ;
         RECT 0.0310 0.1450 0.0530 0.1730 ;
         RECT 0.0310 0.1730 0.0530 0.3000 ;
        RECT 0.0510 0.1310 0.0930 0.1450 ;
         RECT 0.0925 0.1310 0.1145 0.1450 ;
         RECT 0.0925 0.1450 0.1145 0.1730 ;
        RECT 0.0960 0.3190 0.1800 0.3330 ;
        RECT 0.1800 0.0830 0.2610 0.0990 ;
        RECT 0.1800 0.3190 0.2610 0.3330 ;
         RECT 0.2595 0.0830 0.2815 0.0990 ;
         RECT 0.2595 0.0990 0.2815 0.2020 ;
         RECT 0.2595 0.2020 0.2815 0.2300 ;
         RECT 0.2595 0.2300 0.2815 0.3190 ;
         RECT 0.2595 0.3190 0.2815 0.3330 ;
        RECT 0.2800 0.3190 0.6210 0.3330 ;
         RECT 0.6190 0.2020 0.6410 0.2300 ;
         RECT 0.6190 0.2300 0.6410 0.3190 ;
         RECT 0.6190 0.3190 0.6410 0.3330 ;
        RECT 0.6390 0.2020 1.2990 0.2300 ;
        RECT 0.0960 0.2840 0.1380 0.3010 ;
         RECT 0.1360 0.0510 0.1580 0.0650 ;
         RECT 0.1360 0.0650 0.1580 0.1170 ;
         RECT 0.1360 0.1170 0.1580 0.1310 ;
         RECT 0.1360 0.2840 0.1580 0.3010 ;
        RECT 0.1560 0.0510 0.2140 0.0650 ;
        RECT 0.1560 0.1170 0.2140 0.1310 ;
        RECT 0.1560 0.2840 0.2140 0.3010 ;
        RECT 0.2140 0.0510 0.2380 0.0650 ;
        RECT 0.2140 0.1170 0.2380 0.1310 ;
        RECT 0.2140 0.1310 0.2380 0.1360 ;
        RECT 0.2140 0.1360 0.2380 0.1660 ;
        RECT 0.2140 0.1660 0.2380 0.2840 ;
        RECT 0.2140 0.2840 0.2380 0.3010 ;
        RECT 0.2380 0.0510 0.6210 0.0650 ;
         RECT 0.6190 0.0510 0.6410 0.0650 ;
         RECT 0.6190 0.0650 0.6410 0.1170 ;
         RECT 0.6190 0.1170 0.6410 0.1310 ;
         RECT 0.6190 0.1310 0.6410 0.1360 ;
         RECT 0.6190 0.1360 0.6410 0.1660 ;
        RECT 0.6390 0.1360 1.3110 0.1660 ;
      LAYER M1 ;
         RECT 0.0310 0.0360 0.0530 0.1310 ;
         RECT 0.0310 0.1310 0.0530 0.1450 ;
         RECT 0.0310 0.1450 0.0530 0.1730 ;
         RECT 0.0310 0.1730 0.0530 0.3000 ;
        RECT 0.0510 0.1310 0.0930 0.1450 ;
         RECT 0.0925 0.1310 0.1145 0.1450 ;
         RECT 0.0925 0.1450 0.1145 0.1730 ;
        RECT 0.0960 0.3190 0.1800 0.3330 ;
        RECT 0.1800 0.0830 0.2610 0.0990 ;
        RECT 0.1800 0.3190 0.2610 0.3330 ;
         RECT 0.2595 0.0830 0.2815 0.0990 ;
         RECT 0.2595 0.0990 0.2815 0.2020 ;
         RECT 0.2595 0.2020 0.2815 0.2300 ;
         RECT 0.2595 0.2300 0.2815 0.3190 ;
         RECT 0.2595 0.3190 0.2815 0.3330 ;
        RECT 0.2800 0.3190 0.6210 0.3330 ;
         RECT 0.6190 0.2020 0.6410 0.2300 ;
         RECT 0.6190 0.2300 0.6410 0.3190 ;
         RECT 0.6190 0.3190 0.6410 0.3330 ;
        RECT 0.6390 0.2020 1.2990 0.2300 ;
        RECT 0.0960 0.2840 0.1380 0.3010 ;
         RECT 0.1360 0.0510 0.1580 0.0650 ;
         RECT 0.1360 0.0650 0.1580 0.1170 ;
         RECT 0.1360 0.1170 0.1580 0.1310 ;
         RECT 0.1360 0.2840 0.1580 0.3010 ;
        RECT 0.1560 0.0510 0.2140 0.0650 ;
        RECT 0.1560 0.1170 0.2140 0.1310 ;
        RECT 0.1560 0.2840 0.2140 0.3010 ;
        RECT 0.2140 0.0510 0.2380 0.0650 ;
        RECT 0.2140 0.1170 0.2380 0.1310 ;
        RECT 0.2140 0.1310 0.2380 0.1360 ;
        RECT 0.2140 0.1360 0.2380 0.1660 ;
        RECT 0.2140 0.1660 0.2380 0.2840 ;
        RECT 0.2140 0.2840 0.2380 0.3010 ;
        RECT 0.2380 0.0510 0.6210 0.0650 ;
         RECT 0.6190 0.0510 0.6410 0.0650 ;
         RECT 0.6190 0.0650 0.6410 0.1170 ;
         RECT 0.6190 0.1170 0.6410 0.1310 ;
         RECT 0.6190 0.1310 0.6410 0.1360 ;
         RECT 0.6190 0.1360 0.6410 0.1660 ;
        RECT 0.6390 0.1360 1.3110 0.1660 ;
  END
END TBUF_X16

MACRO TIEH
  CLASS core ;
  FOREIGN TIEH 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.1260 BY 0.3840 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0715 0.2360 0.0935 0.3520 ;
         RECT 0.0835 0.2360 0.1055 0.3520 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.0930 0.3980 ;
        RECT 0.0930 0.3700 0.1330 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.1330 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0730 0.0480 0.0950 0.2140 ;
      LAYER M1 ;
         RECT 0.0730 0.0480 0.0950 0.2140 ;
  END
END TIEH

MACRO TIEL
  CLASS core ;
  FOREIGN TIEL 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.1260 BY 0.3840 ;
  PIN Z
    DIRECTION INOUT ;
    PORT
      LAYER M1 ;
        RECT 0.0720 0.0320 0.0960 0.1330 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.0930 0.3980 ;
        RECT 0.0930 0.3700 0.1330 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.1330 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
         RECT 0.0730 0.1680 0.0950 0.3360 ;
      LAYER M1 ;
         RECT 0.0730 0.1680 0.0950 0.3360 ;
  END
END TIEL

MACRO XNOR2_X1
  CLASS core ;
  FOREIGN XNOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.3780 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1165 0.1260 0.1385 0.1400 ;
         RECT 0.1165 0.1400 0.1385 0.2140 ;
        RECT 0.1380 0.1260 0.2430 0.1400 ;
         RECT 0.2410 0.1260 0.2630 0.1400 ;
         RECT 0.2410 0.1400 0.2630 0.2140 ;
         RECT 0.2410 0.2140 0.2630 0.2240 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.1210 0.0530 0.1600 ;
         RECT 0.0310 0.1600 0.0530 0.3380 ;
         RECT 0.0310 0.3380 0.0530 0.3520 ;
        RECT 0.0510 0.3380 0.1800 0.3520 ;
        RECT 0.1800 0.3380 0.3270 0.3520 ;
         RECT 0.3250 0.1600 0.3470 0.3380 ;
         RECT 0.3250 0.3380 0.3470 0.3520 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1790 0.2730 0.2010 0.2740 ;
         RECT 0.1790 0.2740 0.2010 0.3000 ;
         RECT 0.1790 0.3000 0.2010 0.3010 ;
         RECT 0.1975 0.0830 0.2195 0.0970 ;
         RECT 0.1975 0.2730 0.2195 0.2740 ;
         RECT 0.1975 0.2740 0.2195 0.3000 ;
         RECT 0.1975 0.3000 0.2195 0.3010 ;
        RECT 0.2190 0.0830 0.2850 0.0970 ;
        RECT 0.2190 0.2740 0.2850 0.3000 ;
         RECT 0.2830 0.0830 0.3050 0.0970 ;
         RECT 0.2830 0.1240 0.3050 0.1380 ;
         RECT 0.2830 0.1380 0.3050 0.2730 ;
         RECT 0.2830 0.2730 0.3050 0.2740 ;
         RECT 0.2830 0.2740 0.3050 0.3000 ;
         RECT 0.3025 0.0830 0.3245 0.0970 ;
         RECT 0.3025 0.1240 0.3245 0.1380 ;
        RECT 0.3240 0.0830 0.3480 0.0970 ;
        RECT 0.3240 0.0970 0.3480 0.1240 ;
        RECT 0.3240 0.1240 0.3480 0.1380 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.1800 0.3980 ;
        RECT 0.1800 0.3700 0.3510 0.3980 ;
        RECT 0.3510 0.3700 0.3850 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.3850 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.1380 0.0510 0.3510 0.0650 ;
         RECT 0.0730 0.0920 0.0950 0.1080 ;
         RECT 0.0730 0.1080 0.0950 0.1700 ;
         RECT 0.0730 0.1700 0.0950 0.2320 ;
         RECT 0.0730 0.2320 0.0950 0.2460 ;
         RECT 0.0730 0.2460 0.0950 0.2760 ;
        RECT 0.0930 0.0920 0.1540 0.1080 ;
        RECT 0.0930 0.2320 0.1540 0.2460 ;
         RECT 0.1465 0.2320 0.1685 0.2460 ;
         RECT 0.1595 0.1700 0.1815 0.2320 ;
         RECT 0.1595 0.2320 0.1815 0.2460 ;
      LAYER M1 ;
        RECT 0.1380 0.0510 0.3510 0.0650 ;
         RECT 0.0730 0.0920 0.0950 0.1080 ;
         RECT 0.0730 0.1080 0.0950 0.1700 ;
         RECT 0.0730 0.1700 0.0950 0.2320 ;
         RECT 0.0730 0.2320 0.0950 0.2460 ;
         RECT 0.0730 0.2460 0.0950 0.2760 ;
        RECT 0.0930 0.0920 0.1540 0.1080 ;
        RECT 0.0930 0.2320 0.1540 0.2460 ;
         RECT 0.1465 0.2320 0.1685 0.2460 ;
         RECT 0.1595 0.1700 0.1815 0.2320 ;
         RECT 0.1595 0.2320 0.1815 0.2460 ;
  END
END XNOR2_X1

MACRO XOR2_X1
  CLASS core ;
  FOREIGN XOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
  SIZE 0.3780 BY 0.3840 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.1165 0.1720 0.1385 0.2430 ;
         RECT 0.1165 0.2430 0.1385 0.2570 ;
        RECT 0.1380 0.2430 0.1800 0.2570 ;
        RECT 0.1800 0.2430 0.2430 0.2570 ;
         RECT 0.2410 0.1600 0.2630 0.1720 ;
         RECT 0.2410 0.1720 0.2630 0.2430 ;
         RECT 0.2410 0.2430 0.2630 0.2570 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
         RECT 0.0310 0.0320 0.0530 0.0460 ;
         RECT 0.0310 0.0460 0.0530 0.2240 ;
         RECT 0.0310 0.2240 0.0530 0.2630 ;
        RECT 0.0510 0.0320 0.3270 0.0460 ;
         RECT 0.3250 0.0320 0.3470 0.0460 ;
         RECT 0.3250 0.0460 0.3470 0.2240 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1800 0.0820 0.2070 0.1110 ;
         RECT 0.2020 0.0820 0.2240 0.1110 ;
         RECT 0.2020 0.2870 0.2240 0.3010 ;
        RECT 0.2190 0.0820 0.2850 0.1110 ;
        RECT 0.2190 0.2870 0.2850 0.3010 ;
         RECT 0.2830 0.0820 0.3050 0.1110 ;
         RECT 0.2830 0.1110 0.3050 0.2460 ;
         RECT 0.2830 0.2460 0.3050 0.2600 ;
         RECT 0.2830 0.2870 0.3050 0.3010 ;
        RECT 0.3030 0.2460 0.3260 0.2600 ;
        RECT 0.3030 0.2870 0.3260 0.3010 ;
         RECT 0.3250 0.2460 0.3470 0.2600 ;
         RECT 0.3250 0.2600 0.3470 0.2870 ;
         RECT 0.3250 0.2870 0.3470 0.3010 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.3700 0.3510 0.3980 ;
        RECT 0.3510 0.3700 0.3850 0.3980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.0010 0.0010 0.3850 0.0140 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.1610 0.3190 0.3510 0.3330 ;
         RECT 0.0730 0.0680 0.0950 0.1400 ;
         RECT 0.0730 0.1400 0.0950 0.1540 ;
         RECT 0.0730 0.1540 0.0950 0.2160 ;
         RECT 0.0730 0.2160 0.0950 0.2760 ;
         RECT 0.0730 0.2760 0.0950 0.2920 ;
        RECT 0.0930 0.1400 0.1610 0.1540 ;
        RECT 0.0930 0.2760 0.1610 0.2920 ;
         RECT 0.1505 0.1400 0.1725 0.1540 ;
         RECT 0.1505 0.1540 0.1725 0.2160 ;
         RECT 0.1505 0.2760 0.1725 0.2920 ;
         RECT 0.1600 0.1400 0.1820 0.1540 ;
         RECT 0.1600 0.1540 0.1820 0.2160 ;
      LAYER M1 ;
        RECT 0.1610 0.3190 0.3510 0.3330 ;
         RECT 0.0730 0.0680 0.0950 0.1400 ;
         RECT 0.0730 0.1400 0.0950 0.1540 ;
         RECT 0.0730 0.1540 0.0950 0.2160 ;
         RECT 0.0730 0.2160 0.0950 0.2760 ;
         RECT 0.0730 0.2760 0.0950 0.2920 ;
        RECT 0.0930 0.1400 0.1610 0.1540 ;
        RECT 0.0930 0.2760 0.1610 0.2920 ;
         RECT 0.1505 0.1400 0.1725 0.1540 ;
         RECT 0.1505 0.1540 0.1725 0.2160 ;
         RECT 0.1505 0.2760 0.1725 0.2920 ;
         RECT 0.1600 0.1400 0.1820 0.1540 ;
         RECT 0.1600 0.1540 0.1820 0.2160 ;
  END
END XOR2_X1

END LIBRARY
#
# End of file
#
