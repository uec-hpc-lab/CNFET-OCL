VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.001 ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
  LAYER LEF58_PITCH STRING ;
  LAYER LEF58_GAP STRING ;
  LAYER LEF58_EOLKEEPOUT STRING ;
  LAYER LEF58_SPACING STRING ;
  LAYER LEF58_CORNERSPACING STRING ;
  LAYER LEF58_WIDTHTABLE STRING ;
  LAYER LEF58_CUTCLASS STRING ;
  LAYER LEF58_SPACINGTABLE STRING ;
  LAYER LEF58_ENCLOSURE STRING ;
  LAYER LEF58_RIGHTWAYONGRIDONLY STRING ;
  LAYER LEF58_RECTONLY STRING ;
END PROPERTYDEFINITIONS

LAYER nwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE PWELL ;" ;
END pwell


LAYER POLY
  TYPE MASTERSLICE ;
END POLY


LAYER ACT
 TYPE MASTERSLICE ;
END ACT

LAYER V0
TYPE CUT ;
SPACING 0.009 ; 
WIDTH 0.012 ; 
END V0

LAYER M1
  TYPE ROUTING ;
SPACING 0.011 ; 
WIDTH 0.0100 ; 
PITCH 0.021 0.021   ; 
  DIRECTION VERTICAL ;
OFFSET 0.000 0.0105   ; 
END M1

LAYER V1
  TYPE CUT ;
SPACING 0.009 ; 
WIDTH 0.012 ; 

END V1

LAYER MINT1
  TYPE ROUTING ;
SPACING 0.009 ; 
WIDTH 0.012 ; 
PITCH 0.021 0.021   ; 
  DIRECTION HORIZONTAL ;
OFFSET 0.000 0.0105   ; 
END MINT1

LAYER VINT1
  TYPE CUT ;
SPACING 0.009 ; 
WIDTH 0.012 ; 

END VINT1

LAYER MINT2
  TYPE ROUTING ;
SPACING 0.009 ; 
WIDTH 0.012 ; 
PITCH 0.021 0.021   ; 
  DIRECTION VERTICAL ;
OFFSET 0.000 0.0105   ; 
END MINT2

LAYER VINT2
  TYPE CUT ;
SPACING 0.009 ; 
WIDTH 0.012 ; 

END VINT2

LAYER MINT3
  TYPE ROUTING ;
SPACING 0.009 ; 
WIDTH 0.012 ; 
PITCH 0.021 0.021   ; 
  DIRECTION HORIZONTAL ;
OFFSET 0.000 0.0105   ; 
END MINT3

LAYER VINT3
  TYPE CUT ;
SPACING 0.009 ; 
WIDTH 0.012 ; 
END VINT3

LAYER MINT4
  TYPE ROUTING ;
SPACING 0.024 ; 
WIDTH 0.024 ; 
PITCH 0.048 0.048   ; 
  DIRECTION VERTICAL ;
OFFSET 0.000 0.024   ; 
END MINT4

LAYER VINT4
  TYPE CUT ;
SPACING 0.024 ; 
WIDTH 0.024 ; 

END VINT4

LAYER MINT5
  TYPE ROUTING ;
SPACING 0.024 ; 
WIDTH 0.024 ; 
PITCH 0.048 0.048   ; 
  DIRECTION HORIZONTAL ;
OFFSET 0.000 0.024   ; 
END MINT5

LAYER VINT5
  TYPE CUT ;
SPACING 0.024 ; 
WIDTH 0.024 ; 
END VINT5

LAYER MINT6
  TYPE ROUTING ;
SPACING 0.036 ; 
WIDTH 0.036 ; 
PITCH 0.072 0.072   ; 
  DIRECTION  VERTICAL ;
OFFSET 0.000 0.036   ; 
END MINT6

LAYER VINT6
  TYPE CUT ;
SPACING 0.036 ; 
WIDTH 0.036 ; 
END VINT6

LAYER MINT7
  TYPE ROUTING ;
SPACING 0.036 ; 
WIDTH 0.036 ; 
PITCH 0.072 0.072   ; 
  DIRECTION HORIZONTAL ;
OFFSET 0.000 0.036   ; 
END MINT7

LAYER VINT7
  TYPE CUT ;
SPACING 0.036 ; 
WIDTH 0.036 ; 
END VINT7

LAYER MINT8
  TYPE ROUTING ;
SPACING 0.036 ; 
WIDTH 0.036 ; 
PITCH 0.072 0.072  ; 
  DIRECTION VERTICAL ;
OFFSET 0.000 0.036   ; 
END MINT8

VIA V1_0 DEFAULT
  LAYER V1 ;
RECT -0.006 -0.006 0.006 0.006   ; 
  LAYER M1 ;
RECT -0.009 -0.009 0.009 0.009   ; 
  LAYER MINT1 ;
RECT -0.0105 -0.0105 0.0105 0.0105   ; 
END V1_0

VIA VINT1_0 DEFAULT
  LAYER VINT1 ;
RECT -0.006 -0.006 0.006 0.006   ; 
  LAYER MINT1 ;
RECT -0.0105 -0.0105 0.0105 0.0105   ; 
  LAYER MINT2 ;
RECT -0.0105 -0.0105 0.0105 0.0105   ; 
END VINT1_0

VIA VINT2_0 DEFAULT
  LAYER VINT2 ;
RECT -0.006 -0.006 0.006 0.006   ; 
  LAYER MINT2 ;
RECT -0.0105 -0.0105 0.0105 0.0105  ; 
  LAYER MINT3 ;
RECT -0.0105 -0.0105 0.0105 0.0105   ; 
END VINT2_0

VIA VINT3_0 DEFAULT
  LAYER VINT3 ;
RECT -0.006 -0.006 0.006 0.006   ; 
  LAYER MINT3 ;
RECT -0.0105 -0.0105 0.0105 0.0105  ; 
  LAYER MINT4 ;
RECT -0.021 -0.021 0.021 0.021   ; 
END VINT3_0

VIA VINT4_0 DEFAULT
  LAYER VINT4 ;
RECT -0.012 -0.012 0.012 0.012   ; 
  LAYER MINT4 ;
RECT -0.021 -0.021 0.021 0.021   ; 
  LAYER MINT5 ;
RECT -0.021 -0.021 0.021 0.021   ; 
END VINT4_0

VIA VINT5_0 DEFAULT
  LAYER VINT5 ;
RECT -0.012 -0.012 0.012 0.012   ; 
  LAYER MINT5 ;
RECT -0.021 -0.021 0.021 0.021   ; 
  LAYER MINT6 ;
RECT -0.0306 -0.0306 0.0306 0.0306   ; 
END VINT5_0

VIA VINT6_0 DEFAULT
  LAYER VINT6 ;
RECT -0.018 -0.018 0.018 0.018   ; 
  LAYER MINT6 ;
RECT -0.0306 -0.0306 0.0306 0.0306    ; 
  LAYER MINT7 ;
RECT -0.0306 -0.0306 0.0306 0.0306    ; 
END VINT6_0

VIA VINT7_0 DEFAULT
  LAYER VINT7 ;
RECT -0.018 -0.018 0.018 0.018   ; 
  LAYER MINT7 ;
RECT -0.0306 -0.0306 0.0306 0.0306   ; 
  LAYER MINT8 ;
RECT -0.0306 -0.0306 0.0306 0.0306   ; 
END VINT7_0




VIARULE Via1Array-0 GENERATE
  LAYER M1 ;
ENCLOSURE 0.003 0.003   ; 
  LAYER MINT1 ;
ENCLOSURE 0.0015 0.0015   ; 
  LAYER V1 ;
RECT -0.011 -0.011 0.011 0.011   ; 
SPACING 0.010 BY 0.010 ; 
END Via1Array-0

VIARULE Via2Array-0 GENERATE
  LAYER MINT2 ;
ENCLOSURE 0.0045 0.0045   ; 
  LAYER MINT3 ;
ENCLOSURE 0.000 0.000   ; 
  LAYER VINT2 ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.016 BY 0.016 ; 
END Via2Array-0


VIARULE Via3Array-0 GENERATE
  LAYER MINT3 ;
ENCLOSURE 0.0045 0.0045   ; 
  LAYER MINT4 ;
ENCLOSURE 0.0105 0.0105   ; 
  LAYER VINT3 ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.024 BY 0.024 ; 
END Via3Array-0

VIARULE Via4Array-0 GENERATE
  LAYER MINT4 ;
ENCLOSURE 0.009 0.009   ; 
  LAYER MINT5 ;
ENCLOSURE 0.000 0.000   ; 
  LAYER VINT4 ;
RECT -0.012 -0.012 0.012 0.012   ; 
SPACING 0.024 BY 0.024 ; 
END Via4Array-0


VIARULE Via5Array-0 GENERATE
  LAYER MINT5 ;
ENCLOSURE 0.009 0.009   ; 
  LAYER MINT6 ;
ENCLOSURE 0.00906 0.00906   ; 
  LAYER VINT5 ;
RECT -0.012 -0.012 0.012 0.012   ; 
SPACING 0.040 BY 0.040 ; 
END Via5Array-0

VIARULE Via6Array-0 GENERATE
  LAYER MINT6 ;
ENCLOSURE 0.0126 0.0126   ; 
  LAYER MINT7 ;
ENCLOSURE 0.000 0.000   ; 
  LAYER VINT6 ;
RECT -0.020 -0.020 0.020 0.020   ; 
SPACING 0.040 BY 0.040 ; 
END Via6Array-0

VIARULE Via7Array-0 GENERATE
  LAYER MINT7 ;
ENCLOSURE 0.0126 0.0126   ; 
  LAYER MINT8 ;
ENCLOSURE 0.000 0.000   ; 
  LAYER VINT7 ;
RECT -0.020 -0.020 0.020 0.020   ; 
SPACING 0.040 BY 0.040 ; 
END Via7Array-0

VIARULE Via8Array-0 GENERATE
  LAYER MINT1 ;
ENCLOSURE 0.0045 0.0045   ; 
  LAYER MINT2 ;
ENCLOSURE 0.000 0.000   ; 
  LAYER VINT1 ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.016 BY 0.016 ; 
END Via8Array-0


SPACING 
SAMENET M1 M1 0.0105 ; 
SAMENET MINT2 MINT2 0.009 ; 
SAMENET MINT3 MINT3 0.009 ; 
SAMENET MINT4 MINT4 0.024 ; 
SAMENET MINT5 MINT5 0.024 ; 
SAMENET MINT6 MINT6 0.036 ; 
SAMENET MINT7 MINT7 0.036 ; 
SAMENET MINT8 MINT8 0.036 ; 
SAMENET V1 V1 0.009 ; 
SAMENET VINT2 VINT2 0.009 ; 
SAMENET VINT3 VINT3 0.009 ; 
SAMENET VINT4 VINT4 0.024 ; 
SAMENET VINT5 VINT5 0.024 ; 
SAMENET VINT6 VINT6 0.036 ; 
SAMENET VINT7 VINT7 0.036 ; 
SAMENET V1 VINT2 0.000 ; 
SAMENET VINT2 VINT3 0.000 ; 
SAMENET VINT3 VINT4 0.000 ; 
SAMENET VINT4 VINT5 0.000 ; 
SAMENET VINT5 VINT6 0.000 ; 
SAMENET VINT6 VINT7 0.000 ; 
END SPACING



END LIBRARY
#
# End of file
#
