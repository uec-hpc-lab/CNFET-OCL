VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

SITE CORE_TypTyp_0p4_25
  SYMMETRY y ;
  CLASS core ;
SIZE 0.042 BY 0.252 ; 
END CORE_TypTyp_0p4_25



MACRO AND2_X1
  CLASS core ;
  FOREIGN AND2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.084 0.135 0.228   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.041 0.051 0.172   ; 
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.201 0.037 0.219 0.210   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.177 0.261   ; 
RECT 0.177 0.243 0.259 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.259 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.075 0.053 0.093 0.062   ; 
RECT 0.075 0.062 0.093 0.140   ; 
RECT 0.075 0.140 0.093 0.179   ; 
RECT 0.093 0.053 0.159 0.062   ; 
RECT 0.159 0.053 0.177 0.062   ; 
RECT 0.159 0.062 0.177 0.140   ; 
      LAYER M1 ;
RECT 0.075 0.053 0.093 0.062   ; 
RECT 0.075 0.062 0.093 0.140   ; 
RECT 0.075 0.140 0.093 0.179   ; 
RECT 0.093 0.053 0.159 0.062   ; 
RECT 0.159 0.053 0.177 0.062   ; 
RECT 0.159 0.062 0.177 0.140   ; 
  END
END AND2_X1

MACRO AND2_X2
  CLASS core ;
  FOREIGN AND2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.100 0.084 0.116 0.168   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.025 0.081 0.047 0.171   ; 
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.170 0.021 0.172 0.043   ; 
RECT 0.170 0.209 0.172 0.231   ; 
RECT 0.172 0.021 0.188 0.043   ; 
RECT 0.172 0.043 0.188 0.209   ; 
RECT 0.172 0.209 0.188 0.231   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.006 0.243 0.152 0.261   ; 
RECT 0.152 0.243 0.258 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.006 -0.009 0.258 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.030 0.188 0.046 0.198   ; 
RECT 0.046 0.054 0.136 0.064   ; 
RECT 0.046 0.188 0.136 0.198   ; 
RECT 0.136 0.054 0.152 0.064   ; 
RECT 0.136 0.064 0.152 0.188   ; 
RECT 0.136 0.188 0.152 0.198   ; 
      LAYER M1 ;
RECT 0.030 0.188 0.046 0.198   ; 
RECT 0.046 0.054 0.136 0.064   ; 
RECT 0.046 0.188 0.136 0.198   ; 
RECT 0.136 0.054 0.152 0.064   ; 
RECT 0.136 0.064 0.152 0.188   ; 
RECT 0.136 0.188 0.152 0.198   ; 
  END
END AND2_X2


MACRO AND3_X1
  CLASS core ;
  FOREIGN AND3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.336 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.201 0.063 0.219 0.189   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.113 0.063 0.138 0.189   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.032 0.063 0.052 0.189   ; 
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.285 0.037 0.303 0.215   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.261 0.261   ; 
RECT 0.261 0.243 0.343 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.343 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.052 0.033 0.156 0.043   ; 
RECT 0.035 0.207 0.180 0.217   ; 
RECT 0.180 0.032 0.243 0.045   ; 
RECT 0.180 0.207 0.243 0.217   ; 
RECT 0.243 0.032 0.261 0.045   ; 
RECT 0.243 0.045 0.261 0.207   ; 
RECT 0.243 0.207 0.261 0.217   ; 
      LAYER M1 ;
RECT 0.052 0.033 0.156 0.043   ; 
RECT 0.035 0.207 0.180 0.217   ; 
RECT 0.180 0.032 0.243 0.045   ; 
RECT 0.180 0.207 0.243 0.217   ; 
RECT 0.243 0.032 0.261 0.045   ; 
RECT 0.243 0.045 0.261 0.207   ; 
RECT 0.243 0.207 0.261 0.217   ; 
  END
END AND3_X1

MACRO AND3_X2
  CLASS core ;
  FOREIGN AND3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.336 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.105 0.135 0.168   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.030 0.084 0.054 0.168   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.159 0.099 0.177 0.176   ; 
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.240 0.021 0.243 0.051   ; 
RECT 0.240 0.209 0.243 0.231   ; 
RECT 0.243 0.021 0.261 0.051   ; 
RECT 0.243 0.051 0.261 0.209   ; 
RECT 0.243 0.209 0.261 0.231   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.219 0.261   ; 
RECT 0.219 0.243 0.343 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.343 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.032 0.024 0.052 0.051   ; 
RECT 0.032 0.051 0.052 0.062   ; 
RECT 0.052 0.051 0.196 0.062   ; 
RECT 0.035 0.190 0.096 0.201   ; 
RECT 0.096 0.073 0.201 0.083   ; 
RECT 0.096 0.190 0.201 0.201   ; 
RECT 0.201 0.073 0.219 0.083   ; 
RECT 0.201 0.083 0.219 0.190   ; 
RECT 0.201 0.190 0.219 0.201   ; 
      LAYER M1 ;
RECT 0.032 0.024 0.052 0.051   ; 
RECT 0.032 0.051 0.052 0.062   ; 
RECT 0.052 0.051 0.196 0.062   ; 
RECT 0.035 0.190 0.096 0.201   ; 
RECT 0.096 0.073 0.201 0.083   ; 
RECT 0.096 0.190 0.201 0.201   ; 
RECT 0.201 0.073 0.219 0.083   ; 
RECT 0.201 0.083 0.219 0.190   ; 
RECT 0.201 0.190 0.219 0.201   ; 
  END
END AND3_X2

MACRO AND4_X1
  CLASS core ;
  FOREIGN AND4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.378 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.243 0.063 0.261 0.189   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.158 0.063 0.178 0.189   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.063 0.093 0.168   ; 
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.063 0.051 0.189   ; 
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.327 0.037 0.345 0.215   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.303 0.261   ; 
RECT 0.303 0.243 0.385 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.385 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.054 0.209 0.222 0.219   ; 
RECT 0.222 0.033 0.285 0.043   ; 
RECT 0.222 0.209 0.285 0.219   ; 
RECT 0.285 0.033 0.303 0.043   ; 
RECT 0.285 0.043 0.303 0.209   ; 
RECT 0.285 0.209 0.303 0.219   ; 
RECT 0.092 0.033 0.196 0.049   ; 
      LAYER M1 ;
RECT 0.054 0.209 0.222 0.219   ; 
RECT 0.222 0.033 0.285 0.043   ; 
RECT 0.222 0.209 0.285 0.219   ; 
RECT 0.285 0.033 0.303 0.043   ; 
RECT 0.285 0.043 0.303 0.209   ; 
RECT 0.285 0.209 0.303 0.219   ; 
RECT 0.092 0.033 0.196 0.049   ; 
  END
END AND4_X1

MACRO AND4_X2
  CLASS core ;
  FOREIGN AND4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.378 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.219 0.079 0.235 0.189   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.143 0.063 0.159 0.190   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.067 0.063 0.084 0.190   ; 
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.030 0.063 0.046 0.190   ; 
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.294 0.032 0.311 0.210   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.006 0.243 0.273 0.261   ; 
RECT 0.273 0.243 0.384 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.006 -0.009 0.384 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.084 0.033 0.176 0.043   ; 
RECT 0.048 0.209 0.202 0.219   ; 
RECT 0.202 0.054 0.256 0.064   ; 
RECT 0.202 0.209 0.256 0.219   ; 
RECT 0.256 0.054 0.273 0.064   ; 
RECT 0.256 0.064 0.273 0.209   ; 
RECT 0.256 0.209 0.273 0.219   ; 
      LAYER M1 ;
RECT 0.084 0.033 0.176 0.043   ; 
RECT 0.048 0.209 0.202 0.219   ; 
RECT 0.202 0.054 0.256 0.064   ; 
RECT 0.202 0.209 0.256 0.219   ; 
RECT 0.256 0.054 0.273 0.064   ; 
RECT 0.256 0.064 0.273 0.209   ; 
RECT 0.256 0.209 0.273 0.219   ; 
  END
END AND4_X2

MACRO ANTENNA
  CLASS core ;
  FOREIGN ANTENNA 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.126 BY 0.252 ; 
END ANTENNA

MACRO AOI21_X1
  CLASS core ;
  FOREIGN AOI21_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.063 0.135 0.168   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.044 0.051 0.168   ; 
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.201 0.063 0.219 0.168   ; 
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.033 0.093 0.043   ; 
RECT 0.075 0.043 0.093 0.176   ; 
RECT 0.093 0.033 0.201 0.043   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.196 0.261   ; 
RECT 0.196 0.243 0.259 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.259 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.032 0.190 0.052 0.201   ; 
RECT 0.032 0.201 0.052 0.231   ; 
RECT 0.052 0.190 0.196 0.201   ; 
      LAYER M1 ;
RECT 0.032 0.190 0.052 0.201   ; 
RECT 0.032 0.201 0.052 0.231   ; 
RECT 0.052 0.190 0.196 0.201   ; 
  END
END AOI21_X1

MACRO AOI21_X2
  CLASS core ;
  FOREIGN AOI21_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.162 0.099 0.174 0.147   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.106 0.075 0.118 0.085   ; 
RECT 0.106 0.085 0.118 0.147   ; 
RECT 0.106 0.147 0.118 0.168   ; 
RECT 0.118 0.075 0.216 0.085   ; 
RECT 0.216 0.075 0.232 0.085   ; 
RECT 0.216 0.085 0.232 0.147   ; 
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.050 0.084 0.062 0.147   ; 
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.034 0.054 0.078 0.064   ; 
RECT 0.078 0.054 0.090 0.064   ; 
RECT 0.078 0.064 0.090 0.161   ; 
RECT 0.078 0.161 0.090 0.188   ; 
RECT 0.078 0.188 0.090 0.196   ; 
RECT 0.090 0.054 0.188 0.064   ; 
RECT 0.090 0.188 0.188 0.196   ; 
RECT 0.188 0.188 0.190 0.196   ; 
RECT 0.190 0.161 0.202 0.188   ; 
RECT 0.190 0.188 0.202 0.196   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.243 0.230 0.261   ; 
RECT 0.230 0.243 0.234 0.261   ; 
RECT 0.234 0.243 0.256 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.009 0.256 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.021 0.180 0.035 0.209   ; 
RECT 0.021 0.209 0.035 0.219   ; 
RECT 0.035 0.209 0.218 0.219   ; 
RECT 0.218 0.169 0.230 0.180   ; 
RECT 0.218 0.180 0.230 0.209   ; 
RECT 0.218 0.209 0.230 0.219   ; 
RECT 0.064 0.033 0.234 0.043   ; 
      LAYER M1 ;
RECT 0.021 0.180 0.035 0.209   ; 
RECT 0.021 0.209 0.035 0.219   ; 
RECT 0.035 0.209 0.218 0.219   ; 
RECT 0.218 0.169 0.230 0.180   ; 
RECT 0.218 0.180 0.230 0.209   ; 
RECT 0.218 0.209 0.230 0.219   ; 
RECT 0.064 0.033 0.234 0.043   ; 
  END
END AOI21_X2

MACRO AOI22_X1
  CLASS core ;
  FOREIGN AOI22_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.159 0.063 0.177 0.168   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.243 0.063 0.261 0.159   ; 
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.065 0.093 0.189   ; 
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.063 0.051 0.189   ; 
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.092 0.033 0.201 0.043   ; 
RECT 0.201 0.033 0.219 0.043   ; 
RECT 0.201 0.043 0.219 0.191   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.261 0.261   ; 
RECT 0.261 0.243 0.301 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.301 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.054 0.207 0.243 0.221   ; 
RECT 0.243 0.181 0.261 0.207   ; 
RECT 0.243 0.207 0.261 0.221   ; 
      LAYER M1 ;
RECT 0.054 0.207 0.243 0.221   ; 
RECT 0.243 0.181 0.261 0.207   ; 
RECT 0.243 0.207 0.261 0.221   ; 
  END
END AOI22_X1

MACRO AOI22_X2
  CLASS core ;
  FOREIGN AOI22_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.166 0.090 0.177 0.099   ; 
RECT 0.166 0.099 0.177 0.161   ; 
RECT 0.166 0.161 0.177 0.168   ; 
RECT 0.177 0.090 0.250 0.099   ; 
RECT 0.250 0.090 0.264 0.099   ; 
RECT 0.264 0.090 0.275 0.099   ; 
RECT 0.264 0.099 0.275 0.161   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.215 0.121 0.226 0.168   ; 
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.100 0.128 0.173   ; 
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.019 0.079 0.030 0.168   ; 
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.093 0.066 0.103 0.075   ; 
RECT 0.093 0.075 0.103 0.075   ; 
RECT 0.093 0.075 0.103 0.105   ; 
RECT 0.103 0.066 0.139 0.075   ; 
RECT 0.139 0.066 0.142 0.075   ; 
RECT 0.142 0.066 0.152 0.075   ; 
RECT 0.142 0.075 0.152 0.075   ; 
RECT 0.142 0.075 0.152 0.105   ; 
RECT 0.142 0.105 0.152 0.152   ; 
RECT 0.142 0.152 0.152 0.186   ; 
RECT 0.142 0.186 0.152 0.198   ; 
RECT 0.152 0.066 0.240 0.075   ; 
RECT 0.152 0.075 0.240 0.075   ; 
RECT 0.152 0.186 0.240 0.198   ; 
RECT 0.240 0.066 0.250 0.075   ; 
RECT 0.240 0.075 0.250 0.075   ; 
RECT 0.240 0.152 0.250 0.186   ; 
RECT 0.240 0.186 0.250 0.198   ; 
RECT 0.250 0.066 0.264 0.075   ; 
RECT 0.250 0.075 0.264 0.075   ; 
RECT 0.264 0.032 0.275 0.066   ; 
RECT 0.264 0.066 0.275 0.075   ; 
RECT 0.264 0.075 0.275 0.075   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.243 0.275 0.261   ; 
RECT 0.275 0.243 0.298 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.009 0.298 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.155 0.043 0.240 0.054   ; 
RECT 0.240 0.024 0.250 0.043   ; 
RECT 0.240 0.043 0.250 0.054   ; 
RECT 0.029 0.209 0.264 0.219   ; 
RECT 0.264 0.183 0.275 0.209   ; 
RECT 0.264 0.209 0.275 0.219   ; 
RECT 0.033 0.028 0.139 0.047   ; 
      LAYER M1 ;
RECT 0.155 0.043 0.240 0.054   ; 
RECT 0.240 0.024 0.250 0.043   ; 
RECT 0.240 0.043 0.250 0.054   ; 
RECT 0.029 0.209 0.264 0.219   ; 
RECT 0.264 0.183 0.275 0.209   ; 
RECT 0.264 0.209 0.275 0.219   ; 
RECT 0.033 0.028 0.139 0.047   ; 
  END
END AOI22_X2

MACRO BUF_X1
  CLASS core ;
  FOREIGN BUF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.210 BY 0.252 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.063 0.051 0.189   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.158 0.037 0.178 0.231   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.094 0.261   ; 
RECT 0.094 0.243 0.217 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.217 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.075 0.024 0.075 0.060   ; 
RECT 0.075 0.060 0.075 0.070   ; 
RECT 0.075 0.140 0.075 0.150   ; 
RECT 0.075 0.150 0.075 0.183   ; 
RECT 0.075 0.024 0.093 0.060   ; 
RECT 0.075 0.060 0.093 0.070   ; 
RECT 0.075 0.070 0.093 0.140   ; 
RECT 0.075 0.140 0.093 0.150   ; 
RECT 0.075 0.150 0.093 0.183   ; 
RECT 0.093 0.060 0.094 0.070   ; 
RECT 0.093 0.070 0.094 0.140   ; 
RECT 0.093 0.140 0.094 0.150   ; 
      LAYER M1 ;
RECT 0.075 0.024 0.075 0.060   ; 
RECT 0.075 0.060 0.075 0.070   ; 
RECT 0.075 0.140 0.075 0.150   ; 
RECT 0.075 0.150 0.075 0.183   ; 
RECT 0.075 0.024 0.093 0.060   ; 
RECT 0.075 0.060 0.093 0.070   ; 
RECT 0.075 0.070 0.093 0.140   ; 
RECT 0.075 0.140 0.093 0.150   ; 
RECT 0.075 0.150 0.093 0.183   ; 
RECT 0.093 0.060 0.094 0.070   ; 
RECT 0.093 0.070 0.094 0.140   ; 
RECT 0.093 0.140 0.094 0.150   ; 
  END
END BUF_X1

MACRO BUF_X2
  CLASS core ;
  FOREIGN BUF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.210 BY 0.252 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.088 0.051 0.168   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.114 0.198 0.116 0.231   ; 
RECT 0.116 0.024 0.117 0.043   ; 
RECT 0.116 0.198 0.117 0.231   ; 
RECT 0.117 0.024 0.135 0.043   ; 
RECT 0.117 0.043 0.135 0.198   ; 
RECT 0.117 0.198 0.135 0.231   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.093 0.261   ; 
RECT 0.093 0.243 0.217 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.217 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.028 0.182 0.033 0.192   ; 
RECT 0.028 0.192 0.033 0.225   ; 
RECT 0.033 0.032 0.051 0.063   ; 
RECT 0.033 0.063 0.051 0.072   ; 
RECT 0.033 0.182 0.051 0.192   ; 
RECT 0.033 0.192 0.051 0.225   ; 
RECT 0.051 0.063 0.056 0.072   ; 
RECT 0.051 0.182 0.056 0.192   ; 
RECT 0.051 0.192 0.056 0.225   ; 
RECT 0.056 0.063 0.075 0.072   ; 
RECT 0.056 0.182 0.075 0.192   ; 
RECT 0.075 0.063 0.093 0.072   ; 
RECT 0.075 0.072 0.093 0.182   ; 
RECT 0.075 0.182 0.093 0.192   ; 
      LAYER M1 ;
RECT 0.028 0.182 0.033 0.192   ; 
RECT 0.028 0.192 0.033 0.225   ; 
RECT 0.033 0.032 0.051 0.063   ; 
RECT 0.033 0.063 0.051 0.072   ; 
RECT 0.033 0.182 0.051 0.192   ; 
RECT 0.033 0.192 0.051 0.225   ; 
RECT 0.051 0.063 0.056 0.072   ; 
RECT 0.051 0.182 0.056 0.192   ; 
RECT 0.051 0.192 0.056 0.225   ; 
RECT 0.056 0.063 0.075 0.072   ; 
RECT 0.056 0.182 0.075 0.192   ; 
RECT 0.075 0.063 0.093 0.072   ; 
RECT 0.075 0.072 0.093 0.182   ; 
RECT 0.075 0.182 0.093 0.192   ; 
  END
END BUF_X2

MACRO BUF_X4
  CLASS core ;
  FOREIGN BUF_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.210 BY 0.252 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.073 0.079 0.084 0.173   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.059 0.033 0.086 0.043   ; 
RECT 0.086 0.033 0.111 0.043   ; 
RECT 0.086 0.209 0.111 0.219   ; 
RECT 0.111 0.033 0.151 0.043   ; 
RECT 0.111 0.209 0.151 0.219   ; 
RECT 0.151 0.033 0.164 0.043   ; 
RECT 0.151 0.043 0.164 0.209   ; 
RECT 0.151 0.209 0.164 0.219   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.243 0.111 0.261   ; 
RECT 0.111 0.243 0.214 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.009 0.214 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.011 0.054 0.035 0.065   ; 
RECT 0.035 0.054 0.099 0.065   ; 
RECT 0.035 0.187 0.099 0.198   ; 
RECT 0.099 0.054 0.111 0.065   ; 
RECT 0.099 0.065 0.111 0.187   ; 
RECT 0.099 0.187 0.111 0.198   ; 
      LAYER M1 ;
RECT 0.011 0.054 0.035 0.065   ; 
RECT 0.035 0.054 0.099 0.065   ; 
RECT 0.035 0.187 0.099 0.198   ; 
RECT 0.099 0.054 0.111 0.065   ; 
RECT 0.099 0.065 0.111 0.187   ; 
RECT 0.099 0.187 0.111 0.198   ; 
  END
END BUF_X4

MACRO BUF_X8
  CLASS core ;
  FOREIGN BUF_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.210 BY 0.252 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.012 0.084 0.018 0.120   ; 
RECT 0.012 0.120 0.018 0.131   ; 
RECT 0.012 0.131 0.018 0.168   ; 
RECT 0.018 0.120 0.070 0.131   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.079 0.033 0.164 0.043   ; 
RECT 0.079 0.209 0.164 0.219   ; 
RECT 0.164 0.033 0.177 0.043   ; 
RECT 0.164 0.209 0.177 0.219   ; 
RECT 0.177 0.033 0.183 0.043   ; 
RECT 0.177 0.043 0.183 0.209   ; 
RECT 0.177 0.209 0.183 0.219   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 0.243 0.164 0.261   ; 
RECT 0.164 0.243 0.212 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 -0.009 0.212 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.023 0.032 0.027 0.061   ; 
RECT 0.023 0.061 0.027 0.070   ; 
RECT 0.027 0.032 0.033 0.061   ; 
RECT 0.027 0.061 0.033 0.070   ; 
RECT 0.027 0.173 0.033 0.192   ; 
RECT 0.027 0.192 0.033 0.220   ; 
RECT 0.033 0.032 0.037 0.061   ; 
RECT 0.033 0.061 0.037 0.070   ; 
RECT 0.033 0.173 0.037 0.192   ; 
RECT 0.037 0.061 0.083 0.070   ; 
RECT 0.037 0.173 0.083 0.192   ; 
RECT 0.083 0.061 0.090 0.070   ; 
RECT 0.083 0.070 0.090 0.112   ; 
RECT 0.083 0.112 0.090 0.121   ; 
RECT 0.083 0.121 0.090 0.173   ; 
RECT 0.083 0.173 0.090 0.192   ; 
RECT 0.090 0.112 0.164 0.121   ; 
      LAYER M1 ;
RECT 0.023 0.032 0.027 0.061   ; 
RECT 0.023 0.061 0.027 0.070   ; 
RECT 0.027 0.032 0.033 0.061   ; 
RECT 0.027 0.061 0.033 0.070   ; 
RECT 0.027 0.173 0.033 0.192   ; 
RECT 0.027 0.192 0.033 0.220   ; 
RECT 0.033 0.032 0.037 0.061   ; 
RECT 0.033 0.061 0.037 0.070   ; 
RECT 0.033 0.173 0.037 0.192   ; 
RECT 0.037 0.061 0.083 0.070   ; 
RECT 0.037 0.173 0.083 0.192   ; 
RECT 0.083 0.061 0.090 0.070   ; 
RECT 0.083 0.070 0.090 0.112   ; 
RECT 0.083 0.112 0.090 0.121   ; 
RECT 0.083 0.121 0.090 0.173   ; 
RECT 0.083 0.173 0.090 0.192   ; 
RECT 0.090 0.112 0.164 0.121   ; 
  END
END BUF_X8

MACRO BUF_X12
  CLASS core ;
  FOREIGN BUF_X12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.252 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.010 0.077 0.017 0.120   ; 
RECT 0.010 0.120 0.017 0.131   ; 
RECT 0.010 0.131 0.017 0.169   ; 
RECT 0.017 0.120 0.093 0.131   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.102 0.033 0.234 0.043   ; 
RECT 0.102 0.209 0.234 0.219   ; 
RECT 0.234 0.033 0.248 0.043   ; 
RECT 0.234 0.209 0.248 0.219   ; 
RECT 0.248 0.033 0.255 0.043   ; 
RECT 0.248 0.043 0.255 0.209   ; 
RECT 0.248 0.209 0.255 0.219   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 0.243 0.234 0.261   ; 
RECT 0.234 0.243 0.282 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 -0.009 0.282 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.021 0.181 0.024 0.192   ; 
RECT 0.021 0.192 0.024 0.220   ; 
RECT 0.024 0.032 0.031 0.060   ; 
RECT 0.024 0.060 0.031 0.071   ; 
RECT 0.024 0.181 0.031 0.192   ; 
RECT 0.024 0.192 0.031 0.220   ; 
RECT 0.031 0.060 0.034 0.071   ; 
RECT 0.031 0.181 0.034 0.192   ; 
RECT 0.031 0.192 0.034 0.220   ; 
RECT 0.034 0.060 0.101 0.071   ; 
RECT 0.034 0.181 0.101 0.192   ; 
RECT 0.101 0.060 0.107 0.071   ; 
RECT 0.101 0.071 0.107 0.121   ; 
RECT 0.101 0.121 0.107 0.131   ; 
RECT 0.101 0.131 0.107 0.181   ; 
RECT 0.101 0.181 0.107 0.192   ; 
RECT 0.107 0.121 0.234 0.131   ; 
      LAYER M1 ;
RECT 0.021 0.181 0.024 0.192   ; 
RECT 0.021 0.192 0.024 0.220   ; 
RECT 0.024 0.032 0.031 0.060   ; 
RECT 0.024 0.060 0.031 0.071   ; 
RECT 0.024 0.181 0.031 0.192   ; 
RECT 0.024 0.192 0.031 0.220   ; 
RECT 0.031 0.060 0.034 0.071   ; 
RECT 0.031 0.181 0.034 0.192   ; 
RECT 0.031 0.192 0.034 0.220   ; 
RECT 0.034 0.060 0.101 0.071   ; 
RECT 0.034 0.181 0.101 0.192   ; 
RECT 0.101 0.060 0.107 0.071   ; 
RECT 0.101 0.071 0.107 0.121   ; 
RECT 0.101 0.121 0.107 0.131   ; 
RECT 0.101 0.131 0.107 0.181   ; 
RECT 0.101 0.181 0.107 0.192   ; 
RECT 0.107 0.121 0.234 0.131   ; 
  END
END BUF_X12


MACRO BUF_X16
  CLASS core ;
  FOREIGN BUF_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.252 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.008 0.076 0.013 0.117   ; 
RECT 0.008 0.117 0.013 0.135   ; 
RECT 0.008 0.135 0.013 0.168   ; 
RECT 0.013 0.117 0.093 0.135   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.100 0.033 0.245 0.043   ; 
RECT 0.100 0.207 0.245 0.217   ; 
RECT 0.245 0.033 0.256 0.043   ; 
RECT 0.245 0.207 0.256 0.217   ; 
RECT 0.256 0.033 0.261 0.043   ; 
RECT 0.256 0.043 0.261 0.207   ; 
RECT 0.256 0.207 0.261 0.217   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 0.243 0.245 0.261   ; 
RECT 0.245 0.243 0.282 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 -0.009 0.282 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.019 0.032 0.024 0.068   ; 
RECT 0.019 0.068 0.024 0.077   ; 
RECT 0.019 0.150 0.024 0.159   ; 
RECT 0.019 0.159 0.024 0.211   ; 
RECT 0.024 0.068 0.099 0.077   ; 
RECT 0.024 0.150 0.099 0.159   ; 
RECT 0.099 0.068 0.104 0.077   ; 
RECT 0.099 0.077 0.104 0.121   ; 
RECT 0.099 0.121 0.104 0.130   ; 
RECT 0.099 0.130 0.104 0.150   ; 
RECT 0.099 0.150 0.104 0.159   ; 
RECT 0.104 0.121 0.245 0.130   ; 
      LAYER M1 ;
RECT 0.019 0.032 0.024 0.068   ; 
RECT 0.019 0.068 0.024 0.077   ; 
RECT 0.019 0.150 0.024 0.159   ; 
RECT 0.019 0.159 0.024 0.211   ; 
RECT 0.024 0.068 0.099 0.077   ; 
RECT 0.024 0.150 0.099 0.159   ; 
RECT 0.099 0.068 0.104 0.077   ; 
RECT 0.099 0.077 0.104 0.121   ; 
RECT 0.099 0.121 0.104 0.130   ; 
RECT 0.099 0.130 0.104 0.150   ; 
RECT 0.099 0.150 0.104 0.159   ; 
RECT 0.104 0.121 0.245 0.130   ; 
  END
END BUF_X16

MACRO CLKBUF_X1
  CLASS core ;
  FOREIGN CLKBUF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.210 BY 0.252 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.063 0.051 0.189   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.158 0.037 0.178 0.231   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.094 0.261   ; 
RECT 0.094 0.243 0.217 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.217 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.075 0.024 0.075 0.060   ; 
RECT 0.075 0.060 0.075 0.070   ; 
RECT 0.075 0.129 0.075 0.150   ; 
RECT 0.075 0.150 0.075 0.172   ; 
RECT 0.075 0.024 0.093 0.060   ; 
RECT 0.075 0.060 0.093 0.070   ; 
RECT 0.075 0.070 0.093 0.129   ; 
RECT 0.075 0.129 0.093 0.150   ; 
RECT 0.075 0.150 0.093 0.172   ; 
RECT 0.093 0.060 0.094 0.070   ; 
RECT 0.093 0.070 0.094 0.129   ; 
RECT 0.093 0.129 0.094 0.150   ; 
      LAYER M1 ;
RECT 0.075 0.024 0.075 0.060   ; 
RECT 0.075 0.060 0.075 0.070   ; 
RECT 0.075 0.129 0.075 0.150   ; 
RECT 0.075 0.150 0.075 0.172   ; 
RECT 0.075 0.024 0.093 0.060   ; 
RECT 0.075 0.060 0.093 0.070   ; 
RECT 0.075 0.070 0.093 0.129   ; 
RECT 0.075 0.129 0.093 0.150   ; 
RECT 0.075 0.150 0.093 0.172   ; 
RECT 0.093 0.060 0.094 0.070   ; 
RECT 0.093 0.070 0.094 0.129   ; 
RECT 0.093 0.129 0.094 0.150   ; 
  END
END CLKBUF_X1

MACRO CLKBUF_X2
  CLASS core ;
  FOREIGN CLKBUF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.210 BY 0.252 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.097 0.051 0.168   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.114 0.209 0.117 0.231   ; 
RECT 0.117 0.024 0.135 0.209   ; 
RECT 0.117 0.209 0.135 0.231   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.093 0.261   ; 
RECT 0.093 0.243 0.217 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.217 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.032 0.043 0.052 0.063   ; 
RECT 0.032 0.063 0.052 0.072   ; 
RECT 0.032 0.182 0.052 0.192   ; 
RECT 0.032 0.192 0.052 0.225   ; 
RECT 0.052 0.063 0.075 0.072   ; 
RECT 0.052 0.182 0.075 0.192   ; 
RECT 0.075 0.063 0.093 0.072   ; 
RECT 0.075 0.072 0.093 0.182   ; 
RECT 0.075 0.182 0.093 0.192   ; 
      LAYER M1 ;
RECT 0.032 0.043 0.052 0.063   ; 
RECT 0.032 0.063 0.052 0.072   ; 
RECT 0.032 0.182 0.052 0.192   ; 
RECT 0.032 0.192 0.052 0.225   ; 
RECT 0.052 0.063 0.075 0.072   ; 
RECT 0.052 0.182 0.075 0.192   ; 
RECT 0.075 0.063 0.093 0.072   ; 
RECT 0.075 0.072 0.093 0.182   ; 
RECT 0.075 0.182 0.093 0.192   ; 
  END
END CLKBUF_X2

MACRO CLKBUF_X4
  CLASS core ;
  FOREIGN CLKBUF_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.210 BY 0.252 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.047 0.079 0.058 0.173   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.059 0.033 0.084 0.043   ; 
RECT 0.084 0.033 0.084 0.043   ; 
RECT 0.084 0.209 0.084 0.219   ; 
RECT 0.084 0.033 0.151 0.043   ; 
RECT 0.084 0.209 0.151 0.219   ; 
RECT 0.151 0.033 0.164 0.043   ; 
RECT 0.151 0.043 0.164 0.209   ; 
RECT 0.151 0.209 0.164 0.219   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.243 0.084 0.261   ; 
RECT 0.084 0.243 0.214 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.009 0.214 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.017 0.054 0.034 0.064   ; 
RECT 0.034 0.054 0.073 0.064   ; 
RECT 0.034 0.188 0.073 0.198   ; 
RECT 0.073 0.054 0.084 0.064   ; 
RECT 0.073 0.064 0.084 0.188   ; 
RECT 0.073 0.188 0.084 0.198   ; 
      LAYER M1 ;
RECT 0.017 0.054 0.034 0.064   ; 
RECT 0.034 0.054 0.073 0.064   ; 
RECT 0.034 0.188 0.073 0.198   ; 
RECT 0.073 0.054 0.084 0.064   ; 
RECT 0.073 0.064 0.084 0.188   ; 
RECT 0.073 0.188 0.084 0.198   ; 
  END
END CLKBUF_X4

MACRO CLKBUF_X8
  CLASS core ;
  FOREIGN CLKBUF_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.210 BY 0.252 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.012 0.084 0.018 0.108   ; 
RECT 0.012 0.108 0.018 0.117   ; 
RECT 0.012 0.117 0.018 0.168   ; 
RECT 0.018 0.084 0.019 0.108   ; 
RECT 0.018 0.108 0.019 0.117   ; 
RECT 0.019 0.108 0.075 0.117   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.079 0.033 0.168 0.043   ; 
RECT 0.079 0.209 0.168 0.219   ; 
RECT 0.168 0.033 0.177 0.043   ; 
RECT 0.168 0.209 0.177 0.219   ; 
RECT 0.177 0.033 0.183 0.043   ; 
RECT 0.177 0.043 0.183 0.209   ; 
RECT 0.177 0.209 0.183 0.219   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 0.243 0.168 0.261   ; 
RECT 0.168 0.243 0.212 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 -0.009 0.212 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.012 0.054 0.027 0.064   ; 
RECT 0.027 0.054 0.033 0.064   ; 
RECT 0.027 0.148 0.033 0.158   ; 
RECT 0.027 0.158 0.033 0.178   ; 
RECT 0.033 0.054 0.095 0.064   ; 
RECT 0.033 0.148 0.095 0.158   ; 
RECT 0.095 0.054 0.102 0.064   ; 
RECT 0.095 0.064 0.102 0.117   ; 
RECT 0.095 0.117 0.102 0.136   ; 
RECT 0.095 0.136 0.102 0.148   ; 
RECT 0.095 0.148 0.102 0.158   ; 
RECT 0.102 0.117 0.168 0.136   ; 
      LAYER M1 ;
RECT 0.012 0.054 0.027 0.064   ; 
RECT 0.027 0.054 0.033 0.064   ; 
RECT 0.027 0.148 0.033 0.158   ; 
RECT 0.027 0.158 0.033 0.178   ; 
RECT 0.033 0.054 0.095 0.064   ; 
RECT 0.033 0.148 0.095 0.158   ; 
RECT 0.095 0.054 0.102 0.064   ; 
RECT 0.095 0.064 0.102 0.117   ; 
RECT 0.095 0.117 0.102 0.136   ; 
RECT 0.095 0.136 0.102 0.148   ; 
RECT 0.095 0.148 0.102 0.158   ; 
RECT 0.102 0.117 0.168 0.136   ; 
  END
END CLKBUF_X8

MACRO CLKBUF_X12
  CLASS core ;
  FOREIGN CLKBUF_X12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.252 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.010 0.078 0.018 0.110   ; 
RECT 0.010 0.110 0.018 0.121   ; 
RECT 0.010 0.121 0.018 0.174   ; 
RECT 0.018 0.110 0.093 0.121   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.102 0.033 0.218 0.043   ; 
RECT 0.102 0.209 0.218 0.219   ; 
RECT 0.218 0.033 0.248 0.043   ; 
RECT 0.218 0.209 0.248 0.219   ; 
RECT 0.248 0.033 0.255 0.043   ; 
RECT 0.248 0.043 0.255 0.209   ; 
RECT 0.248 0.209 0.255 0.219   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 0.243 0.218 0.261   ; 
RECT 0.218 0.243 0.282 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 -0.009 0.282 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.009 0.054 0.025 0.064   ; 
RECT 0.025 0.054 0.031 0.064   ; 
RECT 0.025 0.180 0.031 0.190   ; 
RECT 0.025 0.190 0.031 0.220   ; 
RECT 0.031 0.054 0.101 0.064   ; 
RECT 0.031 0.180 0.101 0.190   ; 
RECT 0.101 0.054 0.107 0.064   ; 
RECT 0.101 0.064 0.107 0.103   ; 
RECT 0.101 0.103 0.107 0.114   ; 
RECT 0.101 0.114 0.107 0.180   ; 
RECT 0.101 0.180 0.107 0.190   ; 
RECT 0.107 0.054 0.108 0.064   ; 
RECT 0.107 0.064 0.108 0.103   ; 
RECT 0.107 0.103 0.108 0.114   ; 
RECT 0.108 0.103 0.218 0.114   ; 
      LAYER M1 ;
RECT 0.009 0.054 0.025 0.064   ; 
RECT 0.025 0.054 0.031 0.064   ; 
RECT 0.025 0.180 0.031 0.190   ; 
RECT 0.025 0.190 0.031 0.220   ; 
RECT 0.031 0.054 0.101 0.064   ; 
RECT 0.031 0.180 0.101 0.190   ; 
RECT 0.101 0.054 0.107 0.064   ; 
RECT 0.101 0.064 0.107 0.103   ; 
RECT 0.101 0.103 0.107 0.114   ; 
RECT 0.101 0.114 0.107 0.180   ; 
RECT 0.101 0.180 0.107 0.190   ; 
RECT 0.107 0.054 0.108 0.064   ; 
RECT 0.107 0.064 0.108 0.103   ; 
RECT 0.107 0.103 0.108 0.114   ; 
RECT 0.108 0.103 0.218 0.114   ; 
  END
END CLKBUF_X12

MACRO CLKBUF_X16
  CLASS core ;
  FOREIGN CLKBUF_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.252 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.008 0.073 0.013 0.107   ; 
RECT 0.008 0.107 0.013 0.117   ; 
RECT 0.008 0.117 0.013 0.173   ; 
RECT 0.013 0.107 0.093 0.117   ; 
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.100 0.028 0.245 0.047   ; 
RECT 0.100 0.205 0.245 0.224   ; 
RECT 0.245 0.028 0.256 0.047   ; 
RECT 0.245 0.205 0.256 0.224   ; 
RECT 0.256 0.028 0.261 0.047   ; 
RECT 0.256 0.047 0.261 0.205   ; 
RECT 0.256 0.205 0.261 0.224   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 0.243 0.245 0.261   ; 
RECT 0.245 0.243 0.282 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 -0.009 0.282 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.019 0.036 0.024 0.068   ; 
RECT 0.019 0.068 0.024 0.077   ; 
RECT 0.019 0.173 0.024 0.184   ; 
RECT 0.019 0.184 0.024 0.209   ; 
RECT 0.024 0.068 0.100 0.077   ; 
RECT 0.024 0.173 0.100 0.184   ; 
RECT 0.100 0.068 0.110 0.077   ; 
RECT 0.100 0.077 0.110 0.104   ; 
RECT 0.100 0.104 0.110 0.113   ; 
RECT 0.100 0.113 0.110 0.173   ; 
RECT 0.100 0.173 0.110 0.184   ; 
RECT 0.110 0.104 0.245 0.113   ; 
      LAYER M1 ;
RECT 0.019 0.036 0.024 0.068   ; 
RECT 0.019 0.068 0.024 0.077   ; 
RECT 0.019 0.173 0.024 0.184   ; 
RECT 0.019 0.184 0.024 0.209   ; 
RECT 0.024 0.068 0.100 0.077   ; 
RECT 0.024 0.173 0.100 0.184   ; 
RECT 0.100 0.068 0.110 0.077   ; 
RECT 0.100 0.077 0.110 0.104   ; 
RECT 0.100 0.104 0.110 0.113   ; 
RECT 0.100 0.113 0.110 0.173   ; 
RECT 0.100 0.173 0.110 0.184   ; 
RECT 0.110 0.104 0.245 0.113   ; 
  END
END CLKBUF_X16

MACRO DFFRNQ_X1
  CLASS core ;
  FOREIGN DFFRNQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 1.092 BY 0.252 ; 
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.159 0.079 0.177 0.173   ; 
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
RECT 0.462 0.090 0.744 0.099   ; 
RECT 0.744 0.090 0.870 0.099   ; 
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
RECT 0.033 0.084 0.051 0.168   ; 
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 1.040 0.021 1.060 0.231   ; 
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.093 0.261   ; 
RECT 0.093 0.243 0.135 0.261   ; 
RECT 0.135 0.243 0.219 0.261   ; 
RECT 0.219 0.243 0.261 0.261   ; 
RECT 0.261 0.243 0.345 0.261   ; 
RECT 0.345 0.243 0.534 0.261   ; 
RECT 0.534 0.243 0.597 0.261   ; 
RECT 0.597 0.243 0.639 0.261   ; 
RECT 0.639 0.243 0.723 0.261   ; 
RECT 0.723 0.243 0.780 0.261   ; 
RECT 0.780 0.243 0.977 0.261   ; 
RECT 0.977 0.243 1.099 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 1.099 0.009   ; 
    END
  END VSS
  OBS
      LAYER MINT1 ;
RECT 0.096 0.069 0.744 0.078   ; 
RECT 0.054 0.174 0.744 0.183   ; 
      LAYER MINT1 ;
RECT 0.096 0.069 0.744 0.078   ; 
RECT 0.054 0.174 0.744 0.183   ; 
      LAYER M1 ;
RECT 0.117 0.024 0.135 0.228   ; 
RECT 0.201 0.024 0.219 0.228   ; 
RECT 0.348 0.205 0.534 0.223   ; 
RECT 0.285 0.033 0.303 0.043   ; 
RECT 0.285 0.043 0.303 0.144   ; 
RECT 0.285 0.144 0.303 0.220   ; 
RECT 0.303 0.033 0.525 0.043   ; 
RECT 0.525 0.033 0.543 0.043   ; 
RECT 0.525 0.043 0.543 0.144   ; 
RECT 0.378 0.108 0.396 0.166   ; 
RECT 0.378 0.166 0.396 0.175   ; 
RECT 0.396 0.166 0.579 0.175   ; 
RECT 0.579 0.024 0.597 0.108   ; 
RECT 0.579 0.108 0.597 0.166   ; 
RECT 0.579 0.166 0.597 0.175   ; 
RECT 0.579 0.175 0.597 0.221   ; 
RECT 0.663 0.033 0.681 0.043   ; 
RECT 0.663 0.043 0.681 0.120   ; 
RECT 0.663 0.120 0.681 0.220   ; 
RECT 0.681 0.033 0.876 0.043   ; 
RECT 0.876 0.033 0.894 0.043   ; 
RECT 0.876 0.043 0.894 0.120   ; 
RECT 0.803 0.129 0.822 0.209   ; 
RECT 0.803 0.209 0.822 0.219   ; 
RECT 0.822 0.209 0.957 0.219   ; 
RECT 0.957 0.024 0.975 0.043   ; 
RECT 0.957 0.043 0.975 0.129   ; 
RECT 0.957 0.129 0.975 0.209   ; 
RECT 0.957 0.209 0.975 0.219   ; 
RECT 0.975 0.043 0.977 0.129   ; 
RECT 0.975 0.129 0.977 0.209   ; 
RECT 0.975 0.209 0.977 0.219   ; 
RECT 0.032 0.028 0.052 0.046   ; 
RECT 0.032 0.046 0.052 0.055   ; 
RECT 0.032 0.186 0.052 0.199   ; 
RECT 0.032 0.199 0.052 0.225   ; 
RECT 0.052 0.046 0.075 0.055   ; 
RECT 0.052 0.186 0.075 0.199   ; 
RECT 0.075 0.046 0.093 0.055   ; 
RECT 0.075 0.055 0.093 0.186   ; 
RECT 0.075 0.186 0.093 0.199   ; 
RECT 0.243 0.064 0.261 0.162   ; 
RECT 0.327 0.132 0.345 0.188   ; 
RECT 0.345 0.064 0.366 0.096   ; 
RECT 0.483 0.085 0.501 0.144   ; 
RECT 0.621 0.090 0.639 0.190   ; 
RECT 0.705 0.057 0.723 0.104   ; 
RECT 0.705 0.151 0.723 0.204   ; 
RECT 0.759 0.054 0.780 0.225   ; 
RECT 0.831 0.057 0.849 0.104   ; 
      LAYER V1 ;
RECT 0.075 0.174 0.093 0.183   ; 
RECT 0.117 0.069 0.135 0.078   ; 
RECT 0.243 0.069 0.261 0.078   ; 
RECT 0.327 0.174 0.345 0.183   ; 
RECT 0.348 0.069 0.366 0.078   ; 
RECT 0.483 0.090 0.501 0.099   ; 
RECT 0.621 0.174 0.639 0.183   ; 
RECT 0.705 0.069 0.723 0.078   ; 
RECT 0.705 0.174 0.723 0.183   ; 
RECT 0.831 0.090 0.849 0.099   ; 
      LAYER M1 ;
RECT 0.117 0.024 0.135 0.228   ; 
RECT 0.201 0.024 0.219 0.228   ; 
RECT 0.348 0.205 0.534 0.223   ; 
RECT 0.285 0.033 0.303 0.043   ; 
RECT 0.285 0.043 0.303 0.144   ; 
RECT 0.285 0.144 0.303 0.220   ; 
RECT 0.303 0.033 0.525 0.043   ; 
RECT 0.525 0.033 0.543 0.043   ; 
RECT 0.525 0.043 0.543 0.144   ; 
RECT 0.378 0.108 0.396 0.166   ; 
RECT 0.378 0.166 0.396 0.175   ; 
RECT 0.396 0.166 0.579 0.175   ; 
RECT 0.579 0.024 0.597 0.108   ; 
RECT 0.579 0.108 0.597 0.166   ; 
RECT 0.579 0.166 0.597 0.175   ; 
RECT 0.579 0.175 0.597 0.221   ; 
RECT 0.663 0.033 0.681 0.043   ; 
RECT 0.663 0.043 0.681 0.120   ; 
RECT 0.663 0.120 0.681 0.220   ; 
RECT 0.681 0.033 0.876 0.043   ; 
RECT 0.876 0.033 0.894 0.043   ; 
RECT 0.876 0.043 0.894 0.120   ; 
RECT 0.803 0.129 0.822 0.209   ; 
RECT 0.803 0.209 0.822 0.219   ; 
RECT 0.822 0.209 0.957 0.219   ; 
RECT 0.957 0.024 0.975 0.043   ; 
RECT 0.957 0.043 0.975 0.129   ; 
RECT 0.957 0.129 0.975 0.209   ; 
RECT 0.957 0.209 0.975 0.219   ; 
RECT 0.975 0.043 0.977 0.129   ; 
RECT 0.975 0.129 0.977 0.209   ; 
RECT 0.975 0.209 0.977 0.219   ; 
RECT 0.032 0.028 0.052 0.046   ; 
RECT 0.032 0.046 0.052 0.055   ; 
RECT 0.032 0.186 0.052 0.199   ; 
RECT 0.032 0.199 0.052 0.225   ; 
RECT 0.052 0.046 0.075 0.055   ; 
RECT 0.052 0.186 0.075 0.199   ; 
RECT 0.075 0.046 0.093 0.055   ; 
RECT 0.075 0.055 0.093 0.186   ; 
RECT 0.075 0.186 0.093 0.199   ; 
RECT 0.243 0.064 0.261 0.162   ; 
RECT 0.327 0.132 0.345 0.188   ; 
RECT 0.345 0.064 0.366 0.096   ; 
RECT 0.483 0.085 0.501 0.144   ; 
RECT 0.621 0.090 0.639 0.190   ; 
RECT 0.705 0.057 0.723 0.104   ; 
RECT 0.705 0.151 0.723 0.204   ; 
RECT 0.759 0.054 0.780 0.225   ; 
RECT 0.831 0.057 0.849 0.104   ; 
  END
END DFFRNQ_X1

MACRO DFFSNQ_X1
  CLASS core ;
  FOREIGN DFFSNQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 1.092 BY 0.252 ; 
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.159 0.079 0.177 0.173   ; 
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
RECT 0.474 0.090 0.744 0.099   ; 
RECT 0.744 0.090 0.870 0.099   ; 
    END
  END SN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
RECT 0.033 0.084 0.051 0.168   ; 
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 1.040 0.021 1.060 0.231   ; 
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.093 0.261   ; 
RECT 0.093 0.243 0.135 0.261   ; 
RECT 0.135 0.243 0.219 0.261   ; 
RECT 0.219 0.243 0.261 0.261   ; 
RECT 0.261 0.243 0.345 0.261   ; 
RECT 0.345 0.243 0.364 0.261   ; 
RECT 0.364 0.243 0.597 0.261   ; 
RECT 0.597 0.243 0.639 0.261   ; 
RECT 0.639 0.243 0.726 0.261   ; 
RECT 0.726 0.243 0.912 0.261   ; 
RECT 0.912 0.243 0.977 0.261   ; 
RECT 0.977 0.243 1.099 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 1.099 0.009   ; 
    END
  END VSS
  OBS
      LAYER MINT1 ;
RECT 0.096 0.069 0.744 0.078   ; 
RECT 0.054 0.174 0.744 0.183   ; 
      LAYER MINT1 ;
RECT 0.096 0.069 0.744 0.078   ; 
RECT 0.054 0.174 0.744 0.183   ; 
      LAYER M1 ;
RECT 0.117 0.024 0.135 0.228   ; 
RECT 0.201 0.024 0.219 0.228   ; 
RECT 0.285 0.040 0.303 0.049   ; 
RECT 0.285 0.049 0.303 0.120   ; 
RECT 0.285 0.120 0.303 0.220   ; 
RECT 0.303 0.040 0.537 0.049   ; 
RECT 0.537 0.040 0.555 0.049   ; 
RECT 0.537 0.049 0.555 0.120   ; 
RECT 0.621 0.090 0.639 0.188   ; 
RECT 0.705 0.064 0.726 0.106   ; 
RECT 0.705 0.129 0.726 0.195   ; 
RECT 0.831 0.061 0.849 0.104   ; 
RECT 0.789 0.129 0.807 0.188   ; 
RECT 0.789 0.188 0.807 0.198   ; 
RECT 0.807 0.188 0.957 0.198   ; 
RECT 0.957 0.024 0.975 0.043   ; 
RECT 0.957 0.043 0.975 0.129   ; 
RECT 0.957 0.129 0.975 0.188   ; 
RECT 0.957 0.188 0.975 0.198   ; 
RECT 0.975 0.043 0.977 0.129   ; 
RECT 0.975 0.129 0.977 0.188   ; 
RECT 0.975 0.188 0.977 0.198   ; 
RECT 0.030 0.027 0.032 0.045   ; 
RECT 0.030 0.045 0.032 0.058   ; 
RECT 0.032 0.027 0.052 0.045   ; 
RECT 0.032 0.045 0.052 0.058   ; 
RECT 0.032 0.186 0.052 0.199   ; 
RECT 0.032 0.199 0.052 0.225   ; 
RECT 0.052 0.027 0.054 0.045   ; 
RECT 0.052 0.045 0.054 0.058   ; 
RECT 0.052 0.186 0.054 0.199   ; 
RECT 0.054 0.045 0.075 0.058   ; 
RECT 0.054 0.186 0.075 0.199   ; 
RECT 0.075 0.045 0.093 0.058   ; 
RECT 0.075 0.058 0.093 0.186   ; 
RECT 0.075 0.186 0.093 0.199   ; 
RECT 0.243 0.064 0.261 0.162   ; 
RECT 0.327 0.132 0.345 0.194   ; 
RECT 0.345 0.064 0.364 0.100   ; 
RECT 0.495 0.085 0.513 0.120   ; 
RECT 0.399 0.090 0.417 0.188   ; 
RECT 0.399 0.188 0.417 0.198   ; 
RECT 0.417 0.188 0.576 0.198   ; 
RECT 0.576 0.188 0.579 0.198   ; 
RECT 0.576 0.198 0.579 0.225   ; 
RECT 0.579 0.032 0.597 0.090   ; 
RECT 0.579 0.090 0.597 0.188   ; 
RECT 0.579 0.188 0.597 0.198   ; 
RECT 0.579 0.198 0.597 0.225   ; 
RECT 0.663 0.037 0.681 0.047   ; 
RECT 0.663 0.047 0.681 0.120   ; 
RECT 0.663 0.120 0.681 0.221   ; 
RECT 0.681 0.037 0.887 0.047   ; 
RECT 0.887 0.037 0.906 0.047   ; 
RECT 0.887 0.047 0.906 0.120   ; 
RECT 0.726 0.209 0.912 0.219   ; 
      LAYER V1 ;
RECT 0.075 0.174 0.093 0.183   ; 
RECT 0.117 0.069 0.135 0.078   ; 
RECT 0.243 0.069 0.261 0.078   ; 
RECT 0.327 0.174 0.345 0.183   ; 
RECT 0.345 0.069 0.364 0.078   ; 
RECT 0.495 0.090 0.513 0.099   ; 
RECT 0.621 0.174 0.639 0.183   ; 
RECT 0.705 0.069 0.723 0.078   ; 
RECT 0.705 0.174 0.723 0.183   ; 
RECT 0.831 0.090 0.849 0.099   ; 
      LAYER M1 ;
RECT 0.117 0.024 0.135 0.228   ; 
RECT 0.201 0.024 0.219 0.228   ; 
RECT 0.285 0.040 0.303 0.049   ; 
RECT 0.285 0.049 0.303 0.120   ; 
RECT 0.285 0.120 0.303 0.220   ; 
RECT 0.303 0.040 0.537 0.049   ; 
RECT 0.537 0.040 0.555 0.049   ; 
RECT 0.537 0.049 0.555 0.120   ; 
RECT 0.621 0.090 0.639 0.188   ; 
RECT 0.705 0.064 0.726 0.106   ; 
RECT 0.705 0.129 0.726 0.195   ; 
RECT 0.831 0.061 0.849 0.104   ; 
RECT 0.789 0.129 0.807 0.188   ; 
RECT 0.789 0.188 0.807 0.198   ; 
RECT 0.807 0.188 0.957 0.198   ; 
RECT 0.957 0.024 0.975 0.043   ; 
RECT 0.957 0.043 0.975 0.129   ; 
RECT 0.957 0.129 0.975 0.188   ; 
RECT 0.957 0.188 0.975 0.198   ; 
RECT 0.975 0.043 0.977 0.129   ; 
RECT 0.975 0.129 0.977 0.188   ; 
RECT 0.975 0.188 0.977 0.198   ; 
RECT 0.030 0.027 0.032 0.045   ; 
RECT 0.030 0.045 0.032 0.058   ; 
RECT 0.032 0.027 0.052 0.045   ; 
RECT 0.032 0.045 0.052 0.058   ; 
RECT 0.032 0.186 0.052 0.199   ; 
RECT 0.032 0.199 0.052 0.225   ; 
RECT 0.052 0.027 0.054 0.045   ; 
RECT 0.052 0.045 0.054 0.058   ; 
RECT 0.052 0.186 0.054 0.199   ; 
RECT 0.054 0.045 0.075 0.058   ; 
RECT 0.054 0.186 0.075 0.199   ; 
RECT 0.075 0.045 0.093 0.058   ; 
RECT 0.075 0.058 0.093 0.186   ; 
RECT 0.075 0.186 0.093 0.199   ; 
RECT 0.243 0.064 0.261 0.162   ; 
RECT 0.327 0.132 0.345 0.194   ; 
RECT 0.345 0.064 0.364 0.100   ; 
RECT 0.495 0.085 0.513 0.120   ; 
RECT 0.399 0.090 0.417 0.188   ; 
RECT 0.399 0.188 0.417 0.198   ; 
RECT 0.417 0.188 0.576 0.198   ; 
RECT 0.576 0.188 0.579 0.198   ; 
RECT 0.576 0.198 0.579 0.225   ; 
RECT 0.579 0.032 0.597 0.090   ; 
RECT 0.579 0.090 0.597 0.188   ; 
RECT 0.579 0.188 0.597 0.198   ; 
RECT 0.579 0.198 0.597 0.225   ; 
RECT 0.663 0.037 0.681 0.047   ; 
RECT 0.663 0.047 0.681 0.120   ; 
RECT 0.663 0.120 0.681 0.221   ; 
RECT 0.681 0.037 0.887 0.047   ; 
RECT 0.887 0.037 0.906 0.047   ; 
RECT 0.887 0.047 0.906 0.120   ; 
RECT 0.726 0.209 0.912 0.219   ; 
  END
END DFFSNQ_X1

MACRO INV_X1
  CLASS core ;
  FOREIGN INV_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.126 BY 0.252 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.063 0.051 0.189   ; 
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.037 0.093 0.210   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.133 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.133 0.009   ; 
    END
  END VSS
END INV_X1

MACRO INV_X2
  CLASS core ;
  FOREIGN INV_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.126 BY 0.252 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.025 0.063 0.038 0.189   ; 
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.056 0.043 0.070 0.189   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.005 0.243 0.131 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.005 -0.009 0.131 0.009   ; 
    END
  END VSS
END INV_X2

MACRO INV_X4
  CLASS core ;
  FOREIGN INV_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.126 BY 0.252 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.016 0.084 0.026 0.121   ; 
RECT 0.016 0.121 0.026 0.130   ; 
RECT 0.016 0.130 0.026 0.168   ; 
RECT 0.026 0.121 0.078 0.130   ; 
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.013 0.047 0.019 0.066   ; 
RECT 0.019 0.047 0.100 0.066   ; 
RECT 0.019 0.186 0.100 0.205   ; 
RECT 0.100 0.047 0.110 0.066   ; 
RECT 0.100 0.066 0.110 0.186   ; 
RECT 0.100 0.186 0.110 0.205   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.003 0.243 0.129 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.003 -0.009 0.129 0.009   ; 
    END
  END VSS
END INV_X4

MACRO INV_X8
  CLASS core ;
  FOREIGN INV_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.126 BY 0.252 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.022 0.064 0.028 0.130   ; 
RECT 0.022 0.130 0.028 0.150   ; 
RECT 0.022 0.150 0.028 0.189   ; 
RECT 0.028 0.130 0.091 0.150   ; 
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.008 0.207 0.011 0.216   ; 
RECT 0.011 0.036 0.110 0.045   ; 
RECT 0.011 0.207 0.110 0.216   ; 
RECT 0.110 0.036 0.117 0.045   ; 
RECT 0.110 0.045 0.117 0.207   ; 
RECT 0.110 0.207 0.117 0.216   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 0.243 0.128 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 -0.009 0.128 0.009   ; 
    END
  END VSS
END INV_X8

MACRO INV_X12
  CLASS core ;
  FOREIGN INV_X12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.168 BY 0.252 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.021 0.063 0.027 0.121   ; 
RECT 0.021 0.121 0.027 0.130   ; 
RECT 0.021 0.130 0.027 0.189   ; 
RECT 0.027 0.121 0.129 0.130   ; 
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.010 0.033 0.152 0.043   ; 
RECT 0.010 0.209 0.152 0.219   ; 
RECT 0.152 0.033 0.160 0.043   ; 
RECT 0.152 0.043 0.160 0.209   ; 
RECT 0.152 0.209 0.160 0.219   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 0.243 0.170 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.002 -0.009 0.170 0.009   ; 
    END
  END VSS
END INV_X12

MACRO INV_X16
  CLASS core ;
  FOREIGN INV_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.168 BY 0.252 ; 
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.007 0.084 0.011 0.121   ; 
RECT 0.007 0.121 0.011 0.131   ; 
RECT 0.007 0.131 0.011 0.184   ; 
RECT 0.011 0.121 0.137 0.131   ; 
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.001 0.243 0.156 0.261   ; 
RECT 0.156 0.243 0.169 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.001 -0.009 0.169 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.008 0.033 0.151 0.043   ; 
RECT 0.008 0.204 0.151 0.224   ; 
RECT 0.151 0.033 0.156 0.043   ; 
RECT 0.151 0.043 0.156 0.204   ; 
RECT 0.151 0.204 0.156 0.224   ; 
      LAYER M1 ;
RECT 0.008 0.033 0.151 0.043   ; 
RECT 0.008 0.204 0.151 0.224   ; 
RECT 0.151 0.033 0.156 0.043   ; 
RECT 0.151 0.043 0.156 0.204   ; 
RECT 0.151 0.204 0.156 0.224   ; 
  END
END INV_X16

MACRO LHQ_X1
  CLASS core ;
  FOREIGN LHQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.588 BY 0.252 ; 
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.159 0.052 0.177 0.168   ; 
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
RECT 0.033 0.084 0.051 0.168   ; 
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.537 0.043 0.555 0.209   ; 
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.513 0.261   ; 
RECT 0.513 0.243 0.595 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.595 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.032 0.182 0.033 0.192   ; 
RECT 0.032 0.192 0.033 0.231   ; 
RECT 0.033 0.021 0.051 0.030   ; 
RECT 0.033 0.030 0.051 0.060   ; 
RECT 0.033 0.060 0.051 0.070   ; 
RECT 0.033 0.182 0.051 0.192   ; 
RECT 0.033 0.192 0.051 0.231   ; 
RECT 0.051 0.021 0.052 0.030   ; 
RECT 0.051 0.060 0.052 0.070   ; 
RECT 0.051 0.182 0.052 0.192   ; 
RECT 0.051 0.192 0.052 0.231   ; 
RECT 0.052 0.021 0.075 0.030   ; 
RECT 0.052 0.060 0.075 0.070   ; 
RECT 0.052 0.182 0.075 0.192   ; 
RECT 0.075 0.021 0.093 0.030   ; 
RECT 0.075 0.060 0.093 0.070   ; 
RECT 0.075 0.070 0.093 0.106   ; 
RECT 0.075 0.106 0.093 0.115   ; 
RECT 0.075 0.115 0.093 0.136   ; 
RECT 0.075 0.136 0.093 0.182   ; 
RECT 0.075 0.182 0.093 0.192   ; 
RECT 0.093 0.021 0.213 0.030   ; 
RECT 0.213 0.021 0.231 0.030   ; 
RECT 0.213 0.030 0.231 0.060   ; 
RECT 0.213 0.060 0.231 0.070   ; 
RECT 0.213 0.070 0.231 0.106   ; 
RECT 0.213 0.106 0.231 0.115   ; 
RECT 0.231 0.106 0.243 0.115   ; 
RECT 0.243 0.106 0.261 0.115   ; 
RECT 0.243 0.115 0.261 0.136   ; 
RECT 0.348 0.037 0.366 0.047   ; 
RECT 0.348 0.047 0.366 0.162   ; 
RECT 0.366 0.037 0.453 0.047   ; 
RECT 0.453 0.037 0.471 0.047   ; 
RECT 0.453 0.047 0.471 0.162   ; 
RECT 0.453 0.162 0.471 0.194   ; 
RECT 0.117 0.045 0.135 0.151   ; 
RECT 0.117 0.151 0.135 0.182   ; 
RECT 0.117 0.182 0.135 0.192   ; 
RECT 0.135 0.182 0.201 0.192   ; 
RECT 0.201 0.151 0.223 0.182   ; 
RECT 0.201 0.182 0.223 0.192   ; 
RECT 0.180 0.209 0.255 0.219   ; 
RECT 0.255 0.037 0.306 0.056   ; 
RECT 0.255 0.209 0.306 0.219   ; 
RECT 0.306 0.037 0.324 0.056   ; 
RECT 0.306 0.056 0.324 0.100   ; 
RECT 0.306 0.100 0.324 0.209   ; 
RECT 0.306 0.209 0.324 0.209   ; 
RECT 0.306 0.209 0.324 0.219   ; 
RECT 0.324 0.209 0.495 0.209   ; 
RECT 0.324 0.209 0.495 0.219   ; 
RECT 0.495 0.100 0.513 0.209   ; 
RECT 0.495 0.209 0.513 0.209   ; 
RECT 0.495 0.209 0.513 0.219   ; 
      LAYER M1 ;
RECT 0.032 0.182 0.033 0.192   ; 
RECT 0.032 0.192 0.033 0.231   ; 
RECT 0.033 0.021 0.051 0.030   ; 
RECT 0.033 0.030 0.051 0.060   ; 
RECT 0.033 0.060 0.051 0.070   ; 
RECT 0.033 0.182 0.051 0.192   ; 
RECT 0.033 0.192 0.051 0.231   ; 
RECT 0.051 0.021 0.052 0.030   ; 
RECT 0.051 0.060 0.052 0.070   ; 
RECT 0.051 0.182 0.052 0.192   ; 
RECT 0.051 0.192 0.052 0.231   ; 
RECT 0.052 0.021 0.075 0.030   ; 
RECT 0.052 0.060 0.075 0.070   ; 
RECT 0.052 0.182 0.075 0.192   ; 
RECT 0.075 0.021 0.093 0.030   ; 
RECT 0.075 0.060 0.093 0.070   ; 
RECT 0.075 0.070 0.093 0.106   ; 
RECT 0.075 0.106 0.093 0.115   ; 
RECT 0.075 0.115 0.093 0.136   ; 
RECT 0.075 0.136 0.093 0.182   ; 
RECT 0.075 0.182 0.093 0.192   ; 
RECT 0.093 0.021 0.213 0.030   ; 
RECT 0.213 0.021 0.231 0.030   ; 
RECT 0.213 0.030 0.231 0.060   ; 
RECT 0.213 0.060 0.231 0.070   ; 
RECT 0.213 0.070 0.231 0.106   ; 
RECT 0.213 0.106 0.231 0.115   ; 
RECT 0.231 0.106 0.243 0.115   ; 
RECT 0.243 0.106 0.261 0.115   ; 
RECT 0.243 0.115 0.261 0.136   ; 
RECT 0.348 0.037 0.366 0.047   ; 
RECT 0.348 0.047 0.366 0.162   ; 
RECT 0.366 0.037 0.453 0.047   ; 
RECT 0.453 0.037 0.471 0.047   ; 
RECT 0.453 0.047 0.471 0.162   ; 
RECT 0.453 0.162 0.471 0.194   ; 
RECT 0.117 0.045 0.135 0.151   ; 
RECT 0.117 0.151 0.135 0.182   ; 
RECT 0.117 0.182 0.135 0.192   ; 
RECT 0.135 0.182 0.201 0.192   ; 
RECT 0.201 0.151 0.223 0.182   ; 
RECT 0.201 0.182 0.223 0.192   ; 
RECT 0.180 0.209 0.255 0.219   ; 
RECT 0.255 0.037 0.306 0.056   ; 
RECT 0.255 0.209 0.306 0.219   ; 
RECT 0.306 0.037 0.324 0.056   ; 
RECT 0.306 0.056 0.324 0.100   ; 
RECT 0.306 0.100 0.324 0.209   ; 
RECT 0.306 0.209 0.324 0.209   ; 
RECT 0.306 0.209 0.324 0.219   ; 
RECT 0.324 0.209 0.495 0.209   ; 
RECT 0.324 0.209 0.495 0.219   ; 
RECT 0.495 0.100 0.513 0.209   ; 
RECT 0.495 0.209 0.513 0.209   ; 
RECT 0.495 0.209 0.513 0.219   ; 
  END
END LHQ_X1

MACRO MUX2_X1
  CLASS core ;
  FOREIGN MUX2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.546 BY 0.252 ; 
  PIN I0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.369 0.079 0.387 0.173   ; 
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.084 0.093 0.147   ; 
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
RECT 0.077 0.216 0.259 0.225   ; 
      LAYER V1 ;
RECT 0.098 0.216 0.135 0.225   ; 
      LAYER M1 ;
RECT 0.018 0.079 0.036 0.216   ; 
RECT 0.018 0.216 0.036 0.225   ; 
RECT 0.036 0.216 0.146 0.225   ; 
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.453 0.063 0.471 0.209   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.303 0.261   ; 
RECT 0.303 0.243 0.345 0.261   ; 
RECT 0.345 0.243 0.513 0.261   ; 
RECT 0.513 0.243 0.553 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.553 0.009   ; 
    END
  END VSS
  OBS
      LAYER MINT1 ;
RECT 0.180 0.111 0.366 0.120   ; 
      LAYER MINT1 ;
RECT 0.180 0.111 0.366 0.120   ; 
      LAYER M1 ;
RECT 0.052 0.053 0.065 0.062   ; 
RECT 0.065 0.053 0.103 0.062   ; 
RECT 0.065 0.161 0.103 0.171   ; 
RECT 0.065 0.171 0.103 0.189   ; 
RECT 0.103 0.053 0.201 0.062   ; 
RECT 0.103 0.161 0.201 0.171   ; 
RECT 0.201 0.053 0.219 0.062   ; 
RECT 0.201 0.062 0.219 0.161   ; 
RECT 0.201 0.161 0.219 0.171   ; 
RECT 0.190 0.216 0.285 0.231   ; 
RECT 0.285 0.100 0.303 0.216   ; 
RECT 0.285 0.216 0.303 0.231   ; 
RECT 0.327 0.090 0.345 0.140   ; 
RECT 0.243 0.028 0.261 0.048   ; 
RECT 0.243 0.048 0.261 0.162   ; 
RECT 0.243 0.162 0.261 0.201   ; 
RECT 0.261 0.028 0.495 0.048   ; 
RECT 0.495 0.028 0.513 0.048   ; 
RECT 0.495 0.048 0.513 0.162   ; 
      LAYER V1 ;
RECT 0.201 0.111 0.219 0.120   ; 
RECT 0.201 0.216 0.238 0.225   ; 
RECT 0.327 0.111 0.345 0.120   ; 
      LAYER M1 ;
RECT 0.052 0.053 0.065 0.062   ; 
RECT 0.065 0.053 0.103 0.062   ; 
RECT 0.065 0.161 0.103 0.171   ; 
RECT 0.065 0.171 0.103 0.189   ; 
RECT 0.103 0.053 0.201 0.062   ; 
RECT 0.103 0.161 0.201 0.171   ; 
RECT 0.201 0.053 0.219 0.062   ; 
RECT 0.201 0.062 0.219 0.161   ; 
RECT 0.201 0.161 0.219 0.171   ; 
RECT 0.190 0.216 0.285 0.231   ; 
RECT 0.285 0.100 0.303 0.216   ; 
RECT 0.285 0.216 0.303 0.231   ; 
RECT 0.327 0.090 0.345 0.140   ; 
RECT 0.243 0.028 0.261 0.048   ; 
RECT 0.243 0.048 0.261 0.162   ; 
RECT 0.243 0.162 0.261 0.201   ; 
RECT 0.261 0.028 0.495 0.048   ; 
RECT 0.495 0.028 0.513 0.048   ; 
RECT 0.495 0.048 0.513 0.162   ; 
  END
END MUX2_X1

MACRO NAND2_X1
  CLASS core ;
  FOREIGN NAND2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.168 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.084 0.135 0.188   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.084 0.051 0.188   ; 
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.044 0.093 0.063   ; 
RECT 0.075 0.063 0.093 0.209   ; 
RECT 0.093 0.044 0.116 0.063   ; 
RECT 0.116 0.021 0.137 0.044   ; 
RECT 0.116 0.044 0.137 0.063   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.175 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.175 0.009   ; 
    END
  END VSS
END NAND2_X1

MACRO NAND2_X2
  CLASS core ;
  FOREIGN NAND2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.168 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.078 0.074 0.090 0.182   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.022 0.090 0.034 0.222   ; 
RECT 0.022 0.222 0.034 0.231   ; 
RECT 0.034 0.222 0.134 0.231   ; 
RECT 0.134 0.090 0.146 0.222   ; 
RECT 0.134 0.222 0.146 0.231   ; 
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.050 0.041 0.062 0.060   ; 
RECT 0.050 0.060 0.062 0.139   ; 
RECT 0.050 0.139 0.062 0.196   ; 
RECT 0.050 0.196 0.062 0.210   ; 
RECT 0.062 0.041 0.106 0.060   ; 
RECT 0.062 0.196 0.106 0.210   ; 
RECT 0.106 0.041 0.118 0.060   ; 
RECT 0.106 0.139 0.118 0.196   ; 
RECT 0.106 0.196 0.118 0.210   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.243 0.172 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.009 0.172 0.009   ; 
    END
  END VSS
END NAND2_X2

MACRO NAND3_X1
  CLASS core ;
  FOREIGN NAND3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.159 0.105 0.177 0.147   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.084 0.135 0.168   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.071 0.051 0.188   ; 
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.027 0.093 0.036   ; 
RECT 0.075 0.036 0.093 0.084   ; 
RECT 0.075 0.084 0.093 0.168   ; 
RECT 0.075 0.168 0.093 0.222   ; 
RECT 0.075 0.222 0.093 0.231   ; 
RECT 0.093 0.027 0.159 0.036   ; 
RECT 0.093 0.222 0.159 0.231   ; 
RECT 0.159 0.021 0.200 0.027   ; 
RECT 0.159 0.027 0.200 0.036   ; 
RECT 0.159 0.222 0.200 0.231   ; 
RECT 0.200 0.021 0.201 0.027   ; 
RECT 0.200 0.027 0.201 0.036   ; 
RECT 0.200 0.036 0.201 0.084   ; 
RECT 0.200 0.222 0.201 0.231   ; 
RECT 0.201 0.021 0.219 0.027   ; 
RECT 0.201 0.027 0.219 0.036   ; 
RECT 0.201 0.036 0.219 0.084   ; 
RECT 0.201 0.168 0.219 0.222   ; 
RECT 0.201 0.222 0.219 0.231   ; 
RECT 0.219 0.021 0.221 0.027   ; 
RECT 0.219 0.027 0.221 0.036   ; 
RECT 0.219 0.036 0.221 0.084   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.259 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.259 0.009   ; 
    END
  END VSS
END NAND3_X1

MACRO NAND3_X2
  CLASS core ;
  FOREIGN NAND3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.218 0.105 0.230 0.168   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.132 0.081 0.148 0.168   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.050 0.084 0.062 0.168   ; 
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.012 0.186 0.160 0.205   ; 
RECT 0.160 0.186 0.190 0.205   ; 
RECT 0.190 0.061 0.202 0.186   ; 
RECT 0.190 0.186 0.202 0.205   ; 
RECT 0.202 0.186 0.216 0.205   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.243 0.160 0.261   ; 
RECT 0.160 0.243 0.230 0.261   ; 
RECT 0.230 0.243 0.256 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.009 0.256 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.092 0.037 0.218 0.046   ; 
RECT 0.218 0.037 0.230 0.046   ; 
RECT 0.218 0.046 0.230 0.074   ; 
RECT 0.022 0.058 0.160 0.068   ; 
      LAYER M1 ;
RECT 0.092 0.037 0.218 0.046   ; 
RECT 0.218 0.037 0.230 0.046   ; 
RECT 0.218 0.046 0.230 0.074   ; 
RECT 0.022 0.058 0.160 0.068   ; 
  END
END NAND3_X2

MACRO NAND4_X1
  CLASS core ;
  FOREIGN NAND4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.243 0.084 0.261 0.188   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.159 0.079 0.177 0.168   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.064 0.135 0.147   ; 
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.064 0.051 0.188   ; 
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.168 0.093 0.211   ; 
RECT 0.075 0.211 0.093 0.231   ; 
RECT 0.093 0.211 0.201 0.231   ; 
RECT 0.201 0.054 0.219 0.063   ; 
RECT 0.201 0.063 0.219 0.168   ; 
RECT 0.201 0.168 0.219 0.211   ; 
RECT 0.201 0.211 0.219 0.231   ; 
RECT 0.219 0.054 0.240 0.063   ; 
RECT 0.240 0.021 0.264 0.054   ; 
RECT 0.240 0.054 0.264 0.063   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.301 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.301 0.009   ; 
    END
  END VSS
END NAND4_X1

MACRO NAND4_X2
  CLASS core ;
  FOREIGN NAND4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.233 0.117 0.248 0.168   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.155 0.112 0.166 0.173   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.074 0.079 0.086 0.168   ; 
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.021 0.085 0.033 0.168   ; 
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.047 0.182 0.060 0.189   ; 
RECT 0.047 0.189 0.060 0.209   ; 
RECT 0.047 0.209 0.060 0.219   ; 
RECT 0.060 0.209 0.181 0.219   ; 
RECT 0.181 0.096 0.193 0.106   ; 
RECT 0.181 0.106 0.193 0.180   ; 
RECT 0.181 0.180 0.193 0.182   ; 
RECT 0.181 0.182 0.193 0.189   ; 
RECT 0.181 0.209 0.193 0.219   ; 
RECT 0.193 0.096 0.235 0.106   ; 
RECT 0.193 0.180 0.235 0.182   ; 
RECT 0.193 0.182 0.235 0.189   ; 
RECT 0.193 0.209 0.235 0.219   ; 
RECT 0.235 0.096 0.246 0.106   ; 
RECT 0.235 0.180 0.246 0.182   ; 
RECT 0.235 0.182 0.246 0.189   ; 
RECT 0.235 0.189 0.246 0.209   ; 
RECT 0.235 0.209 0.246 0.219   ; 
RECT 0.246 0.096 0.273 0.106   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.243 0.274 0.261   ; 
RECT 0.274 0.243 0.298 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.009 0.298 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.020 0.033 0.033 0.043   ; 
RECT 0.020 0.043 0.033 0.070   ; 
RECT 0.033 0.033 0.180 0.043   ; 
RECT 0.114 0.075 0.261 0.085   ; 
RECT 0.261 0.021 0.274 0.075   ; 
RECT 0.261 0.075 0.274 0.085   ; 
RECT 0.061 0.054 0.206 0.064   ; 
      LAYER M1 ;
RECT 0.020 0.033 0.033 0.043   ; 
RECT 0.020 0.043 0.033 0.070   ; 
RECT 0.033 0.033 0.180 0.043   ; 
RECT 0.114 0.075 0.261 0.085   ; 
RECT 0.261 0.021 0.274 0.075   ; 
RECT 0.261 0.075 0.274 0.085   ; 
RECT 0.061 0.054 0.206 0.064   ; 
  END
END NAND4_X2

MACRO NOR2_X1
  CLASS core ;
  FOREIGN NOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.168 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.064 0.135 0.168   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.064 0.051 0.168   ; 
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.043 0.093 0.189   ; 
RECT 0.075 0.189 0.093 0.209   ; 
RECT 0.093 0.189 0.116 0.209   ; 
RECT 0.116 0.189 0.137 0.209   ; 
RECT 0.116 0.209 0.137 0.231   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.175 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.175 0.009   ; 
    END
  END VSS
END NOR2_X1

MACRO NOR2_X2
  CLASS core ;
  FOREIGN NOR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.168 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.078 0.070 0.090 0.168   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.022 0.021 0.034 0.030   ; 
RECT 0.022 0.030 0.034 0.162   ; 
RECT 0.034 0.021 0.134 0.030   ; 
RECT 0.134 0.021 0.146 0.030   ; 
RECT 0.134 0.030 0.146 0.162   ; 
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.050 0.042 0.062 0.051   ; 
RECT 0.050 0.051 0.062 0.113   ; 
RECT 0.050 0.113 0.062 0.182   ; 
RECT 0.050 0.182 0.062 0.192   ; 
RECT 0.062 0.042 0.077 0.051   ; 
RECT 0.062 0.182 0.077 0.192   ; 
RECT 0.077 0.042 0.091 0.051   ; 
RECT 0.077 0.182 0.091 0.192   ; 
RECT 0.077 0.192 0.091 0.210   ; 
RECT 0.091 0.042 0.106 0.051   ; 
RECT 0.106 0.042 0.118 0.051   ; 
RECT 0.106 0.051 0.118 0.113   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.243 0.172 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.009 0.172 0.009   ; 
    END
  END VSS
END NOR2_X2

MACRO NOR3_X1
  CLASS core ;
  FOREIGN NOR3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.159 0.105 0.177 0.147   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.064 0.135 0.181   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.064 0.051 0.181   ; 
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.021 0.093 0.030   ; 
RECT 0.075 0.030 0.093 0.084   ; 
RECT 0.075 0.084 0.093 0.168   ; 
RECT 0.075 0.168 0.093 0.201   ; 
RECT 0.075 0.201 0.093 0.211   ; 
RECT 0.093 0.021 0.199 0.030   ; 
RECT 0.093 0.201 0.199 0.211   ; 
RECT 0.199 0.021 0.200 0.030   ; 
RECT 0.199 0.030 0.200 0.084   ; 
RECT 0.199 0.201 0.200 0.211   ; 
RECT 0.200 0.021 0.221 0.030   ; 
RECT 0.200 0.030 0.221 0.084   ; 
RECT 0.200 0.168 0.221 0.201   ; 
RECT 0.200 0.201 0.221 0.211   ; 
RECT 0.200 0.211 0.221 0.231   ; 
RECT 0.221 0.021 0.221 0.030   ; 
RECT 0.221 0.030 0.221 0.084   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.259 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.259 0.009   ; 
    END
  END VSS
END NOR3_X1

MACRO NOR3_X2
  CLASS core ;
  FOREIGN NOR3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.218 0.084 0.230 0.147   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.134 0.084 0.146 0.169   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.022 0.084 0.034 0.171   ; 
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.038 0.051 0.190 0.070   ; 
RECT 0.190 0.051 0.202 0.070   ; 
RECT 0.190 0.070 0.202 0.189   ; 
RECT 0.202 0.051 0.214 0.070   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.243 0.230 0.261   ; 
RECT 0.230 0.243 0.256 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.009 0.256 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.092 0.205 0.218 0.215   ; 
RECT 0.218 0.169 0.230 0.205   ; 
RECT 0.218 0.205 0.230 0.215   ; 
RECT 0.038 0.183 0.166 0.194   ; 
      LAYER M1 ;
RECT 0.092 0.205 0.218 0.215   ; 
RECT 0.218 0.169 0.230 0.205   ; 
RECT 0.218 0.205 0.230 0.215   ; 
RECT 0.038 0.183 0.166 0.194   ; 
  END
END NOR3_X2

MACRO NOR4_X1
  CLASS core ;
  FOREIGN NOR4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.243 0.064 0.261 0.168   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.159 0.064 0.177 0.168   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.084 0.135 0.188   ; 
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.064 0.051 0.188   ; 
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.021 0.093 0.033   ; 
RECT 0.075 0.033 0.093 0.071   ; 
RECT 0.093 0.021 0.201 0.033   ; 
RECT 0.201 0.021 0.219 0.033   ; 
RECT 0.201 0.033 0.219 0.071   ; 
RECT 0.201 0.071 0.219 0.189   ; 
RECT 0.201 0.189 0.219 0.198   ; 
RECT 0.219 0.189 0.240 0.198   ; 
RECT 0.240 0.189 0.264 0.198   ; 
RECT 0.240 0.198 0.264 0.231   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.301 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.301 0.009   ; 
    END
  END VSS
END NOR4_X1

MACRO NOR4_X2
  CLASS core ;
  FOREIGN NOR4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.233 0.084 0.248 0.133   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.155 0.079 0.166 0.144   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.101 0.079 0.113 0.173   ; 
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.074 0.084 0.086 0.169   ; 
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.047 0.033 0.060 0.043   ; 
RECT 0.047 0.043 0.060 0.063   ; 
RECT 0.047 0.063 0.060 0.070   ; 
RECT 0.060 0.033 0.181 0.043   ; 
RECT 0.181 0.033 0.193 0.043   ; 
RECT 0.181 0.063 0.193 0.070   ; 
RECT 0.181 0.070 0.193 0.072   ; 
RECT 0.181 0.072 0.193 0.145   ; 
RECT 0.181 0.145 0.193 0.154   ; 
RECT 0.193 0.033 0.235 0.043   ; 
RECT 0.193 0.063 0.235 0.070   ; 
RECT 0.193 0.070 0.235 0.072   ; 
RECT 0.193 0.145 0.235 0.154   ; 
RECT 0.235 0.033 0.246 0.043   ; 
RECT 0.235 0.043 0.246 0.063   ; 
RECT 0.235 0.063 0.246 0.070   ; 
RECT 0.235 0.070 0.246 0.072   ; 
RECT 0.235 0.145 0.246 0.154   ; 
RECT 0.246 0.145 0.277 0.154   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.243 0.180 0.261   ; 
RECT 0.180 0.243 0.206 0.261   ; 
RECT 0.206 0.243 0.274 0.261   ; 
RECT 0.274 0.243 0.298 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.009 0.298 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.088 0.187 0.206 0.198   ; 
RECT 0.020 0.182 0.033 0.209   ; 
RECT 0.020 0.209 0.033 0.219   ; 
RECT 0.033 0.209 0.180 0.219   ; 
RECT 0.141 0.166 0.261 0.175   ; 
RECT 0.261 0.166 0.274 0.175   ; 
RECT 0.261 0.175 0.274 0.225   ; 
      LAYER M1 ;
RECT 0.088 0.187 0.206 0.198   ; 
RECT 0.020 0.182 0.033 0.209   ; 
RECT 0.020 0.209 0.033 0.219   ; 
RECT 0.033 0.209 0.180 0.219   ; 
RECT 0.141 0.166 0.261 0.175   ; 
RECT 0.261 0.166 0.274 0.175   ; 
RECT 0.261 0.175 0.274 0.225   ; 
  END
END NOR4_X2


MACRO OAI21_X1
  CLASS core ;
  FOREIGN OAI21_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.084 0.135 0.189   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.084 0.051 0.208   ; 
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.201 0.084 0.219 0.189   ; 
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.084 0.093 0.209   ; 
RECT 0.075 0.209 0.093 0.219   ; 
RECT 0.093 0.209 0.196 0.219   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.196 0.261   ; 
RECT 0.196 0.243 0.259 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.259 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.033 0.024 0.051 0.051   ; 
RECT 0.033 0.051 0.051 0.062   ; 
RECT 0.051 0.051 0.196 0.062   ; 
      LAYER M1 ;
RECT 0.033 0.024 0.051 0.051   ; 
RECT 0.033 0.051 0.051 0.062   ; 
RECT 0.051 0.051 0.196 0.062   ; 
  END
END OAI21_X1

MACRO OAI21_X2
  CLASS core ;
  FOREIGN OAI21_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.160 0.105 0.176 0.147   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.106 0.079 0.118 0.093   ; 
RECT 0.106 0.093 0.118 0.165   ; 
RECT 0.106 0.165 0.118 0.174   ; 
RECT 0.118 0.165 0.218 0.174   ; 
RECT 0.218 0.093 0.230 0.165   ; 
RECT 0.218 0.165 0.230 0.174   ; 
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.050 0.084 0.062 0.173   ; 
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.013 0.187 0.078 0.198   ; 
RECT 0.078 0.054 0.090 0.064   ; 
RECT 0.078 0.064 0.090 0.091   ; 
RECT 0.078 0.091 0.090 0.187   ; 
RECT 0.078 0.187 0.090 0.198   ; 
RECT 0.090 0.054 0.186 0.064   ; 
RECT 0.090 0.187 0.186 0.198   ; 
RECT 0.186 0.054 0.190 0.064   ; 
RECT 0.190 0.054 0.202 0.064   ; 
RECT 0.190 0.064 0.202 0.091   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.243 0.234 0.261   ; 
RECT 0.234 0.243 0.256 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.009 0.256 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.021 0.033 0.035 0.043   ; 
RECT 0.021 0.043 0.035 0.070   ; 
RECT 0.035 0.033 0.218 0.043   ; 
RECT 0.218 0.033 0.230 0.043   ; 
RECT 0.218 0.043 0.230 0.070   ; 
RECT 0.218 0.070 0.230 0.070   ; 
RECT 0.064 0.209 0.234 0.219   ; 
      LAYER M1 ;
RECT 0.021 0.033 0.035 0.043   ; 
RECT 0.021 0.043 0.035 0.070   ; 
RECT 0.035 0.033 0.218 0.043   ; 
RECT 0.218 0.033 0.230 0.043   ; 
RECT 0.218 0.043 0.230 0.070   ; 
RECT 0.218 0.070 0.230 0.070   ; 
RECT 0.064 0.209 0.234 0.219   ; 
  END
END OAI21_X2

MACRO OAI22_X1
  CLASS core ;
  FOREIGN OAI22_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.159 0.066 0.177 0.189   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.243 0.092 0.261 0.189   ; 
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.063 0.135 0.168   ; 
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.032 0.063 0.052 0.189   ; 
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.092 0.209 0.201 0.219   ; 
RECT 0.201 0.060 0.219 0.209   ; 
RECT 0.201 0.209 0.219 0.219   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.261 0.261   ; 
RECT 0.261 0.243 0.301 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.301 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.033 0.033 0.243 0.043   ; 
RECT 0.243 0.033 0.261 0.043   ; 
RECT 0.243 0.043 0.261 0.070   ; 
      LAYER M1 ;
RECT 0.033 0.033 0.243 0.043   ; 
RECT 0.243 0.033 0.261 0.043   ; 
RECT 0.243 0.043 0.261 0.070   ; 
  END
END OAI22_X1

MACRO OAI22_X2
  CLASS core ;
  FOREIGN OAI22_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.166 0.084 0.177 0.091   ; 
RECT 0.166 0.091 0.177 0.153   ; 
RECT 0.166 0.153 0.177 0.162   ; 
RECT 0.177 0.153 0.264 0.162   ; 
RECT 0.264 0.091 0.275 0.153   ; 
RECT 0.264 0.153 0.275 0.162   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.215 0.084 0.226 0.131   ; 
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.079 0.128 0.159   ; 
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.044 0.079 0.054 0.168   ; 
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.093 0.127 0.103 0.174   ; 
RECT 0.093 0.174 0.103 0.183   ; 
RECT 0.103 0.174 0.142 0.183   ; 
RECT 0.142 0.056 0.152 0.064   ; 
RECT 0.142 0.064 0.152 0.091   ; 
RECT 0.142 0.091 0.152 0.127   ; 
RECT 0.142 0.127 0.152 0.174   ; 
RECT 0.142 0.174 0.152 0.183   ; 
RECT 0.152 0.056 0.240 0.064   ; 
RECT 0.152 0.174 0.240 0.183   ; 
RECT 0.240 0.056 0.250 0.064   ; 
RECT 0.240 0.064 0.250 0.091   ; 
RECT 0.240 0.174 0.250 0.183   ; 
RECT 0.250 0.174 0.264 0.183   ; 
RECT 0.264 0.174 0.275 0.183   ; 
RECT 0.264 0.183 0.275 0.221   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 0.243 0.139 0.261   ; 
RECT 0.139 0.243 0.250 0.261   ; 
RECT 0.250 0.243 0.275 0.261   ; 
RECT 0.275 0.243 0.298 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.004 -0.009 0.298 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.154 0.198 0.240 0.209   ; 
RECT 0.240 0.198 0.250 0.209   ; 
RECT 0.240 0.209 0.250 0.228   ; 
RECT 0.016 0.033 0.264 0.043   ; 
RECT 0.264 0.033 0.275 0.043   ; 
RECT 0.264 0.043 0.275 0.069   ; 
RECT 0.019 0.201 0.139 0.220   ; 
      LAYER M1 ;
RECT 0.154 0.198 0.240 0.209   ; 
RECT 0.240 0.198 0.250 0.209   ; 
RECT 0.240 0.209 0.250 0.228   ; 
RECT 0.016 0.033 0.264 0.043   ; 
RECT 0.264 0.033 0.275 0.043   ; 
RECT 0.264 0.043 0.275 0.069   ; 
RECT 0.019 0.201 0.139 0.220   ; 
  END
END OAI22_X2

MACRO OR2_X1
  CLASS core ;
  FOREIGN OR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.032 0.135 0.168   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.080 0.051 0.210   ; 
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.201 0.037 0.219 0.210   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.177 0.261   ; 
RECT 0.177 0.243 0.259 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.259 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.075 0.043 0.093 0.110   ; 
RECT 0.075 0.110 0.093 0.182   ; 
RECT 0.075 0.182 0.093 0.192   ; 
RECT 0.093 0.182 0.159 0.192   ; 
RECT 0.159 0.110 0.177 0.182   ; 
RECT 0.159 0.182 0.177 0.192   ; 
      LAYER M1 ;
RECT 0.075 0.043 0.093 0.110   ; 
RECT 0.075 0.110 0.093 0.182   ; 
RECT 0.075 0.182 0.093 0.192   ; 
RECT 0.093 0.182 0.159 0.192   ; 
RECT 0.159 0.110 0.177 0.182   ; 
RECT 0.159 0.182 0.177 0.192   ; 
  END
END OR2_X1

MACRO OR2_X2
  CLASS core ;
  FOREIGN OR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.064 0.079 0.080 0.168   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.028 0.084 0.044 0.168   ; 
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.170 0.021 0.172 0.045   ; 
RECT 0.170 0.209 0.172 0.231   ; 
RECT 0.172 0.021 0.188 0.045   ; 
RECT 0.172 0.045 0.188 0.209   ; 
RECT 0.172 0.209 0.188 0.231   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.006 0.243 0.152 0.261   ; 
RECT 0.152 0.243 0.258 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.006 -0.009 0.258 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.043 0.051 0.082 0.062   ; 
RECT 0.082 0.051 0.136 0.062   ; 
RECT 0.082 0.190 0.136 0.199   ; 
RECT 0.136 0.051 0.152 0.062   ; 
RECT 0.136 0.062 0.152 0.190   ; 
RECT 0.136 0.190 0.152 0.199   ; 
      LAYER M1 ;
RECT 0.043 0.051 0.082 0.062   ; 
RECT 0.082 0.051 0.136 0.062   ; 
RECT 0.082 0.190 0.136 0.199   ; 
RECT 0.136 0.051 0.152 0.062   ; 
RECT 0.136 0.062 0.152 0.190   ; 
RECT 0.136 0.190 0.152 0.199   ; 
  END
END OR2_X2

MACRO OR3_X1
  CLASS core ;
  FOREIGN OR3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.336 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.201 0.063 0.219 0.189   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.116 0.063 0.137 0.189   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.030 0.063 0.054 0.189   ; 
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.285 0.037 0.303 0.215   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.154 0.261   ; 
RECT 0.154 0.243 0.261 0.261   ; 
RECT 0.261 0.243 0.343 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.343 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.035 0.036 0.182 0.045   ; 
RECT 0.182 0.036 0.243 0.045   ; 
RECT 0.182 0.207 0.243 0.221   ; 
RECT 0.243 0.036 0.261 0.045   ; 
RECT 0.243 0.045 0.261 0.207   ; 
RECT 0.243 0.207 0.261 0.221   ; 
RECT 0.056 0.209 0.154 0.219   ; 
      LAYER M1 ;
RECT 0.035 0.036 0.182 0.045   ; 
RECT 0.182 0.036 0.243 0.045   ; 
RECT 0.182 0.207 0.243 0.221   ; 
RECT 0.243 0.036 0.261 0.045   ; 
RECT 0.243 0.045 0.261 0.207   ; 
RECT 0.243 0.207 0.261 0.221   ; 
RECT 0.056 0.209 0.154 0.219   ; 
  END
END OR3_X1

MACRO OR3_X2
  CLASS core ;
  FOREIGN OR3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.336 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.084 0.093 0.147   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.084 0.051 0.173   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.159 0.076 0.177 0.147   ; 
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.240 0.021 0.243 0.043   ; 
RECT 0.240 0.209 0.243 0.231   ; 
RECT 0.243 0.021 0.261 0.043   ; 
RECT 0.243 0.043 0.261 0.209   ; 
RECT 0.243 0.209 0.261 0.231   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.198 0.261   ; 
RECT 0.198 0.243 0.219 0.261   ; 
RECT 0.219 0.243 0.343 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.343 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.033 0.188 0.051 0.198   ; 
RECT 0.033 0.198 0.051 0.225   ; 
RECT 0.051 0.188 0.198 0.198   ; 
RECT 0.039 0.051 0.092 0.062   ; 
RECT 0.092 0.051 0.201 0.062   ; 
RECT 0.092 0.165 0.201 0.176   ; 
RECT 0.201 0.051 0.219 0.062   ; 
RECT 0.201 0.062 0.219 0.165   ; 
RECT 0.201 0.165 0.219 0.176   ; 
      LAYER M1 ;
RECT 0.033 0.188 0.051 0.198   ; 
RECT 0.033 0.198 0.051 0.225   ; 
RECT 0.051 0.188 0.198 0.198   ; 
RECT 0.039 0.051 0.092 0.062   ; 
RECT 0.092 0.051 0.201 0.062   ; 
RECT 0.092 0.165 0.201 0.176   ; 
RECT 0.201 0.051 0.219 0.062   ; 
RECT 0.201 0.062 0.219 0.165   ; 
RECT 0.201 0.165 0.219 0.176   ; 
  END
END OR3_X2

MACRO OR4_X1
  CLASS core ;
  FOREIGN OR4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.378 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.243 0.063 0.261 0.189   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.158 0.063 0.178 0.189   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.075 0.065 0.093 0.189   ; 
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.063 0.051 0.189   ; 
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.327 0.037 0.345 0.210   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.196 0.261   ; 
RECT 0.196 0.243 0.303 0.261   ; 
RECT 0.303 0.243 0.385 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.385 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.035 0.033 0.222 0.043   ; 
RECT 0.222 0.033 0.285 0.043   ; 
RECT 0.222 0.207 0.285 0.217   ; 
RECT 0.285 0.033 0.303 0.043   ; 
RECT 0.285 0.043 0.303 0.207   ; 
RECT 0.285 0.207 0.303 0.217   ; 
RECT 0.096 0.202 0.196 0.215   ; 
      LAYER M1 ;
RECT 0.035 0.033 0.222 0.043   ; 
RECT 0.222 0.033 0.285 0.043   ; 
RECT 0.222 0.207 0.285 0.217   ; 
RECT 0.285 0.033 0.303 0.043   ; 
RECT 0.285 0.043 0.303 0.207   ; 
RECT 0.285 0.207 0.303 0.217   ; 
RECT 0.096 0.202 0.196 0.215   ; 
  END
END OR4_X1

MACRO OR4_X2
  CLASS core ;
  FOREIGN OR4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.378 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.181 0.063 0.197 0.174   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.143 0.070 0.159 0.189   ; 
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.067 0.070 0.084 0.189   ; 
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.030 0.062 0.046 0.189   ; 
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.293 0.042 0.312 0.231   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.006 0.243 0.178 0.261   ; 
RECT 0.178 0.243 0.272 0.261   ; 
RECT 0.272 0.243 0.384 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.006 -0.009 0.384 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.086 0.205 0.178 0.224   ; 
RECT 0.032 0.028 0.202 0.047   ; 
RECT 0.202 0.028 0.255 0.047   ; 
RECT 0.202 0.186 0.255 0.205   ; 
RECT 0.255 0.028 0.272 0.047   ; 
RECT 0.255 0.047 0.272 0.186   ; 
RECT 0.255 0.186 0.272 0.205   ; 
      LAYER M1 ;
RECT 0.086 0.205 0.178 0.224   ; 
RECT 0.032 0.028 0.202 0.047   ; 
RECT 0.202 0.028 0.255 0.047   ; 
RECT 0.202 0.186 0.255 0.205   ; 
RECT 0.255 0.028 0.272 0.047   ; 
RECT 0.255 0.047 0.272 0.186   ; 
RECT 0.255 0.186 0.272 0.205   ; 
  END
END OR4_X2



MACRO TIEH
  CLASS core ;
  FOREIGN TIEH 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.126 BY 0.252 ; 
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.072 0.155 0.093 0.231   ; 
RECT 0.093 0.155 0.096 0.231   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.093 0.261   ; 
RECT 0.093 0.243 0.133 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.133 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.075 0.032 0.093 0.140   ; 
      LAYER M1 ;
RECT 0.075 0.032 0.093 0.140   ; 
  END
END TIEH

MACRO TIEL
  CLASS core ;
  FOREIGN TIEL 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.126 BY 0.252 ; 
  PIN Z
    DIRECTION INOUT ;
    PORT
      LAYER M1 ;
RECT 0.072 0.021 0.096 0.087   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.093 0.261   ; 
RECT 0.093 0.243 0.133 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.133 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.075 0.110 0.093 0.221   ; 
      LAYER M1 ;
RECT 0.075 0.110 0.093 0.221   ; 
  END
END TIEL

MACRO XNOR2_X1
  CLASS core ;
  FOREIGN XNOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.378 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.083 0.138 0.092   ; 
RECT 0.117 0.092 0.138 0.140   ; 
RECT 0.138 0.083 0.243 0.092   ; 
RECT 0.243 0.083 0.261 0.092   ; 
RECT 0.243 0.092 0.261 0.140   ; 
RECT 0.243 0.140 0.261 0.147   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.079 0.051 0.105   ; 
RECT 0.033 0.105 0.051 0.222   ; 
RECT 0.033 0.222 0.051 0.231   ; 
RECT 0.051 0.222 0.180 0.231   ; 
RECT 0.180 0.222 0.327 0.231   ; 
RECT 0.327 0.105 0.345 0.222   ; 
RECT 0.327 0.222 0.345 0.231   ; 
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.182 0.179 0.198 0.180   ; 
RECT 0.182 0.180 0.198 0.197   ; 
RECT 0.182 0.197 0.198 0.198   ; 
RECT 0.198 0.054 0.219 0.064   ; 
RECT 0.198 0.179 0.219 0.180   ; 
RECT 0.198 0.180 0.219 0.197   ; 
RECT 0.198 0.197 0.219 0.198   ; 
RECT 0.219 0.054 0.285 0.064   ; 
RECT 0.219 0.180 0.285 0.197   ; 
RECT 0.285 0.054 0.303 0.064   ; 
RECT 0.285 0.081 0.303 0.091   ; 
RECT 0.285 0.091 0.303 0.179   ; 
RECT 0.285 0.179 0.303 0.180   ; 
RECT 0.285 0.180 0.303 0.197   ; 
RECT 0.303 0.054 0.324 0.064   ; 
RECT 0.303 0.081 0.324 0.091   ; 
RECT 0.324 0.054 0.348 0.064   ; 
RECT 0.324 0.064 0.348 0.081   ; 
RECT 0.324 0.081 0.348 0.091   ; 
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.180 0.261   ; 
RECT 0.180 0.243 0.351 0.261   ; 
RECT 0.351 0.243 0.385 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.385 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.138 0.033 0.351 0.043   ; 
RECT 0.075 0.060 0.093 0.071   ; 
RECT 0.075 0.071 0.093 0.112   ; 
RECT 0.075 0.112 0.093 0.152   ; 
RECT 0.075 0.152 0.093 0.161   ; 
RECT 0.075 0.161 0.093 0.181   ; 
RECT 0.093 0.060 0.154 0.071   ; 
RECT 0.093 0.152 0.154 0.161   ; 
RECT 0.154 0.152 0.161 0.161   ; 
RECT 0.161 0.112 0.180 0.152   ; 
RECT 0.161 0.152 0.180 0.161   ; 
      LAYER M1 ;
RECT 0.138 0.033 0.351 0.043   ; 
RECT 0.075 0.060 0.093 0.071   ; 
RECT 0.075 0.071 0.093 0.112   ; 
RECT 0.075 0.112 0.093 0.152   ; 
RECT 0.075 0.152 0.093 0.161   ; 
RECT 0.075 0.161 0.093 0.181   ; 
RECT 0.093 0.060 0.154 0.071   ; 
RECT 0.093 0.152 0.154 0.161   ; 
RECT 0.154 0.152 0.161 0.161   ; 
RECT 0.161 0.112 0.180 0.152   ; 
RECT 0.161 0.152 0.180 0.161   ; 
  END
END XNOR2_X1

MACRO XOR2_X1
  CLASS core ;
  FOREIGN XOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.378 BY 0.252 ; 
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.117 0.113 0.138 0.159   ; 
RECT 0.117 0.159 0.138 0.169   ; 
RECT 0.138 0.159 0.180 0.169   ; 
RECT 0.180 0.159 0.243 0.169   ; 
RECT 0.243 0.105 0.261 0.113   ; 
RECT 0.243 0.113 0.261 0.159   ; 
RECT 0.243 0.159 0.261 0.169   ; 
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
RECT 0.033 0.021 0.051 0.030   ; 
RECT 0.033 0.030 0.051 0.147   ; 
RECT 0.033 0.147 0.051 0.173   ; 
RECT 0.051 0.021 0.327 0.030   ; 
RECT 0.327 0.021 0.345 0.030   ; 
RECT 0.327 0.030 0.345 0.147   ; 
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
RECT 0.180 0.054 0.207 0.054   ; 
RECT 0.180 0.054 0.207 0.073   ; 
RECT 0.207 0.054 0.219 0.054   ; 
RECT 0.207 0.054 0.219 0.073   ; 
RECT 0.207 0.188 0.219 0.198   ; 
RECT 0.219 0.054 0.285 0.073   ; 
RECT 0.219 0.188 0.285 0.198   ; 
RECT 0.285 0.054 0.303 0.073   ; 
RECT 0.285 0.073 0.303 0.161   ; 
RECT 0.285 0.161 0.303 0.171   ; 
RECT 0.285 0.188 0.303 0.198   ; 
RECT 0.303 0.161 0.326 0.171   ; 
RECT 0.303 0.188 0.326 0.198   ; 
RECT 0.326 0.161 0.346 0.171   ; 
RECT 0.326 0.171 0.346 0.188   ; 
RECT 0.326 0.188 0.346 0.198   ; 
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 0.243 0.351 0.261   ; 
RECT 0.351 0.243 0.385 0.261   ; 
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
RECT -0.007 -0.009 0.385 0.009   ; 
    END
  END VSS
  OBS
      LAYER M1 ;
RECT 0.161 0.209 0.351 0.219   ; 
RECT 0.075 0.045 0.093 0.092   ; 
RECT 0.075 0.092 0.093 0.101   ; 
RECT 0.075 0.101 0.093 0.142   ; 
RECT 0.075 0.142 0.093 0.181   ; 
RECT 0.075 0.181 0.093 0.192   ; 
RECT 0.093 0.092 0.161 0.101   ; 
RECT 0.093 0.181 0.161 0.192   ; 
RECT 0.161 0.092 0.162 0.101   ; 
RECT 0.161 0.101 0.162 0.142   ; 
RECT 0.161 0.181 0.162 0.192   ; 
RECT 0.162 0.092 0.180 0.101   ; 
RECT 0.162 0.101 0.180 0.142   ; 
      LAYER M1 ;
RECT 0.161 0.209 0.351 0.219   ; 
RECT 0.075 0.045 0.093 0.092   ; 
RECT 0.075 0.092 0.093 0.101   ; 
RECT 0.075 0.101 0.093 0.142   ; 
RECT 0.075 0.142 0.093 0.181   ; 
RECT 0.075 0.181 0.093 0.192   ; 
RECT 0.093 0.092 0.161 0.101   ; 
RECT 0.093 0.181 0.161 0.192   ; 
RECT 0.161 0.092 0.162 0.101   ; 
RECT 0.161 0.101 0.162 0.142   ; 
RECT 0.161 0.181 0.162 0.192   ; 
RECT 0.162 0.092 0.180 0.101   ; 
RECT 0.162 0.101 0.180 0.142   ; 
  END
END XOR2_X1

END LIBRARY
#
# End of file
#
