# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2014, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *       NGLibraryCreator, Development_version_64 - build 201405300513        *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on us19.nangate.us for user Lucio Rech (lre).
# Local time is now Tue, 3 Jun 2014, 13:07:07.
# Main process id is 12480.

VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

SITE CORE_TypTyp_0p4_25
  SYMMETRY y ;
  CLASS core ;
SIZE 0.042 BY 0.504 ;
END CORE_TypTyp_0p4_25

MACRO AND2_X1
  CLASS core ;
  FOREIGN AND2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.168 0.135187 0.456685 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.0833435 0.0511875 0.34453 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.200812 0.0748125 0.219187 0.42 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.177187 0.522375 ;
  RECT 0.177187 0.485625 0.258562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.258562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0748125 0.106312 0.093122 0.124687 ;
  RECT 0.0748125 0.124687 0.093122 0.280875 ;
  RECT 0.0748125 0.280875 0.093122 0.357 ;
  RECT 0.093122 0.106312 0.158812 0.124687 ;
  RECT 0.158812 0.106312 0.177187 0.124687 ;
  RECT 0.158812 0.124687 0.177187 0.280875 ;
      LAYER M1 ;
  RECT 0.0748125 0.106312 0.093122 0.124687 ;
  RECT 0.0748125 0.124687 0.093122 0.280875 ;
  RECT 0.0748125 0.280875 0.093122 0.357 ;
  RECT 0.093122 0.106312 0.158812 0.124687 ;
  RECT 0.158812 0.106312 0.177187 0.124687 ;
  RECT 0.158812 0.124687 0.177187 0.280875 ;
  END
END AND2_X1

MACRO AND2_X2
  CLASS core ;
  FOREIGN AND2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.168 0.135187 0.336 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0295312 0.16275 0.054469 0.34125 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.198187 0.042 0.200812 0.0853125 ;
  RECT 0.198187 0.418687 0.200812 0.462 ;
  RECT 0.200812 0.042 0.219187 0.0853125 ;
  RECT 0.200812 0.0853125 0.219187 0.418687 ;
  RECT 0.200812 0.418687 0.219187 0.462 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.177187 0.522375 ;
  RECT 0.177187 0.485625 0.300563 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.300563 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0354375 0.376688 0.0538125 0.395062 ;
  RECT 0.0538125 0.108937 0.158812 0.127312 ;
  RECT 0.0538125 0.376688 0.158812 0.395062 ;
  RECT 0.158812 0.108937 0.177187 0.127312 ;
  RECT 0.158812 0.127312 0.177187 0.376688 ;
  RECT 0.158812 0.376688 0.177187 0.395062 ;
      LAYER M1 ;
  RECT 0.0354375 0.376688 0.0538125 0.395062 ;
  RECT 0.0538125 0.108937 0.158812 0.127312 ;
  RECT 0.0538125 0.376688 0.158812 0.395062 ;
  RECT 0.158812 0.108937 0.177187 0.127312 ;
  RECT 0.158812 0.127312 0.177187 0.376688 ;
  RECT 0.158812 0.376688 0.177187 0.395062 ;
  END
END AND2_X2

MACRO AND3_X1
  CLASS core ;
  FOREIGN AND3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.336 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.200812 0.126 0.219187 0.378 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.113466 0.126 0.138469 0.378 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0315 0.126 0.0525 0.378 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.284813 0.0748125 0.303187 0.429187 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.261188 0.522375 ;
  RECT 0.261188 0.485625 0.342562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.342562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.051844 0.065625 0.156187 0.086625 ;
  RECT 0.0354375 0.414095 0.179812 0.43247 ;
  RECT 0.179812 0.062344 0.242812 0.089906 ;
  RECT 0.179812 0.414095 0.242812 0.43247 ;
  RECT 0.242812 0.062344 0.261188 0.089906 ;
  RECT 0.242812 0.089906 0.261188 0.414095 ;
  RECT 0.242812 0.414095 0.261188 0.43247 ;
      LAYER M1 ;
  RECT 0.051844 0.065625 0.156187 0.086625 ;
  RECT 0.0354375 0.414095 0.179812 0.43247 ;
  RECT 0.179812 0.062344 0.242812 0.089906 ;
  RECT 0.179812 0.414095 0.242812 0.43247 ;
  RECT 0.242812 0.062344 0.261188 0.089906 ;
  RECT 0.242812 0.089906 0.261188 0.414095 ;
  RECT 0.242812 0.414095 0.261188 0.43247 ;
  END
END AND3_X1

MACRO AND3_X2
  CLASS core ;
  FOREIGN AND3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.336 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.21 0.135187 0.336655 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0295312 0.168 0.054469 0.336 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.198187 0.177187 0.352405 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.240187 0.042 0.242812 0.103031 ;
  RECT 0.240187 0.418687 0.242812 0.462 ;
  RECT 0.242812 0.042 0.261188 0.103031 ;
  RECT 0.242812 0.103031 0.261188 0.418687 ;
  RECT 0.242812 0.418687 0.261188 0.462 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.219187 0.522375 ;
  RECT 0.219187 0.485625 0.342562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.342562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0315 0.04725 0.0525 0.102375 ;
  RECT 0.0315 0.102375 0.0525 0.123375 ;
  RECT 0.0525 0.102375 0.195562 0.123375 ;
  RECT 0.0354375 0.38128 0.0958125 0.40228 ;
  RECT 0.0958125 0.147 0.200812 0.165375 ;
  RECT 0.0958125 0.38128 0.200812 0.40228 ;
  RECT 0.200812 0.147 0.219187 0.165375 ;
  RECT 0.200812 0.165375 0.219187 0.38128 ;
  RECT 0.200812 0.38128 0.219187 0.40228 ;
      LAYER M1 ;
  RECT 0.0315 0.04725 0.0525 0.102375 ;
  RECT 0.0315 0.102375 0.0525 0.123375 ;
  RECT 0.0525 0.102375 0.195562 0.123375 ;
  RECT 0.0354375 0.38128 0.0958125 0.40228 ;
  RECT 0.0958125 0.147 0.200812 0.165375 ;
  RECT 0.0958125 0.38128 0.200812 0.40228 ;
  RECT 0.200812 0.147 0.219187 0.165375 ;
  RECT 0.200812 0.165375 0.219187 0.38128 ;
  RECT 0.200812 0.38128 0.219187 0.40228 ;
  END
END AND3_X2

MACRO AND4_X1
  CLASS core ;
  FOREIGN AND4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.378 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.242812 0.126 0.261188 0.378 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.1575 0.126 0.1785 0.378 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.126 0.093122 0.336 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.126 0.0511875 0.378 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.326813 0.0748125 0.345187 0.429187 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.303187 0.522375 ;
  RECT 0.303187 0.485625 0.384562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.384562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0538125 0.417375 0.221812 0.438375 ;
  RECT 0.221812 0.065625 0.284813 0.086625 ;
  RECT 0.221812 0.417375 0.284813 0.438375 ;
  RECT 0.284813 0.065625 0.303187 0.086625 ;
  RECT 0.284813 0.086625 0.303187 0.417375 ;
  RECT 0.284813 0.417375 0.303187 0.438375 ;
  RECT 0.0924655 0.064969 0.195562 0.096469 ;
      LAYER M1 ;
  RECT 0.0538125 0.417375 0.221812 0.438375 ;
  RECT 0.221812 0.065625 0.284813 0.086625 ;
  RECT 0.221812 0.417375 0.284813 0.438375 ;
  RECT 0.284813 0.065625 0.303187 0.086625 ;
  RECT 0.284813 0.086625 0.303187 0.417375 ;
  RECT 0.284813 0.417375 0.303187 0.438375 ;
  RECT 0.0924655 0.064969 0.195562 0.096469 ;
  END
END AND4_X1

MACRO AND4_X2
  CLASS core ;
  FOREIGN AND4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.42 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.242812 0.158156 0.261188 0.378 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.126 0.177187 0.378655 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.126 0.093122 0.378655 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.126 0.0511875 0.378655 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.326813 0.063 0.345187 0.42 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.303187 0.522375 ;
  RECT 0.303187 0.485625 0.426563 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.426563 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.093122 0.065625 0.195562 0.086625 ;
  RECT 0.0538125 0.417375 0.224437 0.438375 ;
  RECT 0.224437 0.108281 0.284813 0.129281 ;
  RECT 0.224437 0.417375 0.284813 0.438375 ;
  RECT 0.284813 0.108281 0.303187 0.129281 ;
  RECT 0.284813 0.129281 0.303187 0.417375 ;
  RECT 0.284813 0.417375 0.303187 0.438375 ;
      LAYER M1 ;
  RECT 0.093122 0.065625 0.195562 0.086625 ;
  RECT 0.0538125 0.417375 0.224437 0.438375 ;
  RECT 0.224437 0.108281 0.284813 0.129281 ;
  RECT 0.224437 0.417375 0.284813 0.438375 ;
  RECT 0.284813 0.108281 0.303187 0.129281 ;
  RECT 0.284813 0.129281 0.303187 0.417375 ;
  RECT 0.284813 0.417375 0.303187 0.438375 ;
  END
END AND4_X2

MACRO ANTENNA
  CLASS core ;
  FOREIGN ANTENNA 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.126 BY 0.504 ;
END ANTENNA

MACRO AOI21_X1
  CLASS core ;
  FOREIGN AOI21_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.126 0.135187 0.336 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.0879375 0.0511875 0.336 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.200812 0.126 0.219187 0.336 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.065625 0.093122 0.086625 ;
  RECT 0.0748125 0.086625 0.093122 0.35175 ;
  RECT 0.093122 0.065625 0.200812 0.086625 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.195562 0.522375 ;
  RECT 0.195562 0.485625 0.258562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.258562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0315 0.380625 0.0525 0.401625 ;
  RECT 0.0315 0.401625 0.0525 0.462 ;
  RECT 0.0525 0.380625 0.195562 0.401625 ;
      LAYER M1 ;
  RECT 0.0315 0.380625 0.0525 0.401625 ;
  RECT 0.0315 0.401625 0.0525 0.462 ;
  RECT 0.0525 0.380625 0.195562 0.401625 ;
  END
END AOI21_X1

MACRO AOI21_X2
  CLASS core ;
  FOREIGN AOI21_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.378 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.242812 0.198187 0.261188 0.294 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.150937 0.177187 0.169312 ;
  RECT 0.158812 0.169312 0.177187 0.294 ;
  RECT 0.158812 0.294 0.177187 0.336 ;
  RECT 0.177187 0.150937 0.32353 0.169312 ;
  RECT 0.32353 0.150937 0.34847 0.169312 ;
  RECT 0.32353 0.169312 0.34847 0.294 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.168 0.093122 0.294 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.050531 0.108937 0.116812 0.127312 ;
  RECT 0.116812 0.108937 0.135187 0.127312 ;
  RECT 0.116812 0.127312 0.135187 0.320905 ;
  RECT 0.116812 0.320905 0.135187 0.374652 ;
  RECT 0.116812 0.374652 0.135187 0.393095 ;
  RECT 0.135187 0.108937 0.282187 0.127312 ;
  RECT 0.135187 0.374652 0.282187 0.393095 ;
  RECT 0.282187 0.374652 0.284813 0.393095 ;
  RECT 0.284813 0.320905 0.303187 0.374652 ;
  RECT 0.284813 0.374652 0.303187 0.393095 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.345187 0.522375 ;
  RECT 0.345187 0.485625 0.351095 0.522375 ;
  RECT 0.351095 0.485625 0.384562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.384562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0315 0.360938 0.0525 0.41672 ;
  RECT 0.0315 0.41672 0.0525 0.43903 ;
  RECT 0.0525 0.41672 0.326813 0.43903 ;
  RECT 0.326813 0.338625 0.345187 0.360938 ;
  RECT 0.326813 0.360938 0.345187 0.41672 ;
  RECT 0.326813 0.41672 0.345187 0.43903 ;
  RECT 0.0958125 0.066872 0.351095 0.0853125 ;
      LAYER M1 ;
  RECT 0.0315 0.360938 0.0525 0.41672 ;
  RECT 0.0315 0.41672 0.0525 0.43903 ;
  RECT 0.0525 0.41672 0.326813 0.43903 ;
  RECT 0.326813 0.338625 0.345187 0.360938 ;
  RECT 0.326813 0.360938 0.345187 0.41672 ;
  RECT 0.326813 0.41672 0.345187 0.43903 ;
  RECT 0.0958125 0.066872 0.351095 0.0853125 ;
  END
END AOI21_X2

MACRO AOI22_X1
  CLASS core ;
  FOREIGN AOI22_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.126 0.177187 0.336 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.242812 0.126 0.261188 0.31828 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.129937 0.093122 0.378 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.126 0.0511875 0.378 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0924655 0.066872 0.200812 0.0853125 ;
  RECT 0.200812 0.066872 0.219187 0.0853125 ;
  RECT 0.200812 0.0853125 0.219187 0.381937 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.261188 0.522375 ;
  RECT 0.261188 0.485625 0.300563 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.300563 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0538125 0.413438 0.242812 0.442312 ;
  RECT 0.242812 0.362905 0.261188 0.413438 ;
  RECT 0.242812 0.413438 0.261188 0.442312 ;
      LAYER M1 ;
  RECT 0.0538125 0.413438 0.242812 0.442312 ;
  RECT 0.242812 0.362905 0.261188 0.413438 ;
  RECT 0.242812 0.413438 0.261188 0.442312 ;
  END
END AOI22_X1

MACRO AOI22_X2
  CLASS core ;
  FOREIGN AOI22_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.504 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.284813 0.179812 0.303187 0.198187 ;
  RECT 0.284813 0.198187 0.303187 0.320905 ;
  RECT 0.284813 0.320905 0.303187 0.336 ;
  RECT 0.303187 0.179812 0.429187 0.198187 ;
  RECT 0.429187 0.179812 0.452748 0.198187 ;
  RECT 0.452748 0.179812 0.471187 0.198187 ;
  RECT 0.452748 0.198187 0.471187 0.320905 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.368812 0.242812 0.387188 0.336 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.200812 0.200812 0.219187 0.345187 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.158812 0.0511875 0.336 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.13125 0.177187 0.149625 ;
  RECT 0.158812 0.149625 0.177187 0.150281 ;
  RECT 0.158812 0.150281 0.177187 0.21 ;
  RECT 0.177187 0.13125 0.237562 0.149625 ;
  RECT 0.237562 0.13125 0.242812 0.149625 ;
  RECT 0.242812 0.13125 0.261188 0.149625 ;
  RECT 0.242812 0.149625 0.261188 0.150281 ;
  RECT 0.242812 0.150281 0.261188 0.21 ;
  RECT 0.242812 0.21 0.261188 0.303845 ;
  RECT 0.242812 0.303845 0.261188 0.372685 ;
  RECT 0.242812 0.372685 0.261188 0.395062 ;
  RECT 0.261188 0.13125 0.410813 0.149625 ;
  RECT 0.261188 0.149625 0.410813 0.150281 ;
  RECT 0.261188 0.372685 0.410813 0.395062 ;
  RECT 0.410813 0.13125 0.429187 0.149625 ;
  RECT 0.410813 0.149625 0.429187 0.150281 ;
  RECT 0.410813 0.303845 0.429187 0.372685 ;
  RECT 0.410813 0.372685 0.429187 0.395062 ;
  RECT 0.429187 0.13125 0.452748 0.149625 ;
  RECT 0.429187 0.149625 0.452748 0.150281 ;
  RECT 0.452748 0.063 0.471187 0.13125 ;
  RECT 0.452748 0.13125 0.471187 0.149625 ;
  RECT 0.452748 0.149625 0.471187 0.150281 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.471187 0.522375 ;
  RECT 0.471187 0.485625 0.510565 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.510565 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.266437 0.086625 0.410813 0.107625 ;
  RECT 0.410813 0.04725 0.429187 0.086625 ;
  RECT 0.410813 0.086625 0.429187 0.107625 ;
  RECT 0.050531 0.418687 0.452748 0.437063 ;
  RECT 0.452748 0.36553 0.471187 0.418687 ;
  RECT 0.452748 0.418687 0.471187 0.437063 ;
  RECT 0.056372 0.057028 0.237562 0.095156 ;
      LAYER M1 ;
  RECT 0.266437 0.086625 0.410813 0.107625 ;
  RECT 0.410813 0.04725 0.429187 0.086625 ;
  RECT 0.410813 0.086625 0.429187 0.107625 ;
  RECT 0.050531 0.418687 0.452748 0.437063 ;
  RECT 0.452748 0.36553 0.471187 0.418687 ;
  RECT 0.452748 0.418687 0.471187 0.437063 ;
  RECT 0.056372 0.057028 0.237562 0.095156 ;
  END
END AOI22_X2

MACRO BUF_X1
  CLASS core ;
  FOREIGN BUF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.21 BY 0.504 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.126 0.0511875 0.378 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.1575 0.0748125 0.1785 0.462 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.093778 0.522375 ;
  RECT 0.093778 0.485625 0.216562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.216562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0748125 0.04725 0.075469 0.121406 ;
  RECT 0.0748125 0.121406 0.075469 0.139781 ;
  RECT 0.0748125 0.280875 0.075469 0.29925 ;
  RECT 0.0748125 0.29925 0.075469 0.366187 ;
  RECT 0.075469 0.04725 0.093122 0.121406 ;
  RECT 0.075469 0.121406 0.093122 0.139781 ;
  RECT 0.075469 0.139781 0.093122 0.280875 ;
  RECT 0.075469 0.280875 0.093122 0.29925 ;
  RECT 0.075469 0.29925 0.093122 0.366187 ;
  RECT 0.093122 0.121406 0.093778 0.139781 ;
  RECT 0.093122 0.139781 0.093778 0.280875 ;
  RECT 0.093122 0.280875 0.093778 0.29925 ;
      LAYER M1 ;
  RECT 0.0748125 0.04725 0.075469 0.121406 ;
  RECT 0.0748125 0.121406 0.075469 0.139781 ;
  RECT 0.0748125 0.280875 0.075469 0.29925 ;
  RECT 0.0748125 0.29925 0.075469 0.366187 ;
  RECT 0.075469 0.04725 0.093122 0.121406 ;
  RECT 0.075469 0.121406 0.093122 0.139781 ;
  RECT 0.075469 0.139781 0.093122 0.280875 ;
  RECT 0.075469 0.280875 0.093122 0.29925 ;
  RECT 0.075469 0.29925 0.093122 0.366187 ;
  RECT 0.093122 0.121406 0.093778 0.139781 ;
  RECT 0.093122 0.139781 0.093778 0.280875 ;
  RECT 0.093122 0.280875 0.093778 0.29925 ;
  END
END BUF_X1

MACRO BUF_X2
  CLASS core ;
  FOREIGN BUF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.21 BY 0.504 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.175219 0.0511875 0.336 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.114122 0.39572 0.116156 0.462 ;
  RECT 0.116156 0.04725 0.116812 0.086625 ;
  RECT 0.116156 0.39572 0.116812 0.462 ;
  RECT 0.116812 0.04725 0.135187 0.086625 ;
  RECT 0.116812 0.086625 0.135187 0.39572 ;
  RECT 0.116812 0.39572 0.135187 0.462 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.093122 0.522375 ;
  RECT 0.093122 0.485625 0.216562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.216562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0275625 0.364875 0.0328125 0.38325 ;
  RECT 0.0275625 0.38325 0.0328125 0.450188 ;
  RECT 0.0328125 0.063 0.0511875 0.126 ;
  RECT 0.0328125 0.126 0.0511875 0.144375 ;
  RECT 0.0328125 0.364875 0.0511875 0.38325 ;
  RECT 0.0328125 0.38325 0.0511875 0.450188 ;
  RECT 0.0511875 0.126 0.056372 0.144375 ;
  RECT 0.0511875 0.364875 0.056372 0.38325 ;
  RECT 0.0511875 0.38325 0.056372 0.450188 ;
  RECT 0.056372 0.126 0.0748125 0.144375 ;
  RECT 0.056372 0.364875 0.0748125 0.38325 ;
  RECT 0.0748125 0.126 0.093122 0.144375 ;
  RECT 0.0748125 0.144375 0.093122 0.364875 ;
  RECT 0.0748125 0.364875 0.093122 0.38325 ;
      LAYER M1 ;
  RECT 0.0275625 0.364875 0.0328125 0.38325 ;
  RECT 0.0275625 0.38325 0.0328125 0.450188 ;
  RECT 0.0328125 0.063 0.0511875 0.126 ;
  RECT 0.0328125 0.126 0.0511875 0.144375 ;
  RECT 0.0328125 0.364875 0.0511875 0.38325 ;
  RECT 0.0328125 0.38325 0.0511875 0.450188 ;
  RECT 0.0511875 0.126 0.056372 0.144375 ;
  RECT 0.0511875 0.364875 0.056372 0.38325 ;
  RECT 0.0511875 0.38325 0.056372 0.450188 ;
  RECT 0.056372 0.126 0.0748125 0.144375 ;
  RECT 0.056372 0.364875 0.0748125 0.38325 ;
  RECT 0.0748125 0.126 0.093122 0.144375 ;
  RECT 0.0748125 0.144375 0.093122 0.364875 ;
  RECT 0.0748125 0.364875 0.093122 0.38325 ;
  END
END BUF_X2

MACRO BUF_X4
  CLASS core ;
  FOREIGN BUF_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.336 BY 0.504 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.158812 0.135187 0.345187 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.095156 0.066872 0.137812 0.0853125 ;
  RECT 0.137812 0.066872 0.177187 0.0853125 ;
  RECT 0.137812 0.418687 0.177187 0.437063 ;
  RECT 0.177187 0.066872 0.2415 0.0853125 ;
  RECT 0.177187 0.418687 0.2415 0.437063 ;
  RECT 0.2415 0.066872 0.2625 0.0853125 ;
  RECT 0.2415 0.0853125 0.2625 0.418687 ;
  RECT 0.2415 0.418687 0.2625 0.437063 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.177187 0.522375 ;
  RECT 0.177187 0.485625 0.342562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.342562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0177187 0.108937 0.056372 0.129937 ;
  RECT 0.056372 0.108937 0.158812 0.129937 ;
  RECT 0.056372 0.373997 0.158812 0.395062 ;
  RECT 0.158812 0.108937 0.177187 0.129937 ;
  RECT 0.158812 0.129937 0.177187 0.373997 ;
  RECT 0.158812 0.373997 0.177187 0.395062 ;
      LAYER M1 ;
  RECT 0.0177187 0.108937 0.056372 0.129937 ;
  RECT 0.056372 0.108937 0.158812 0.129937 ;
  RECT 0.056372 0.373997 0.158812 0.395062 ;
  RECT 0.158812 0.108937 0.177187 0.129937 ;
  RECT 0.158812 0.129937 0.177187 0.373997 ;
  RECT 0.158812 0.373997 0.177187 0.395062 ;
  END
END BUF_X4

MACRO BUF_X8
  CLASS core ;
  FOREIGN BUF_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.588 BY 0.504 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.168 0.0511875 0.240187 ;
  RECT 0.0328125 0.240187 0.0511875 0.261188 ;
  RECT 0.0328125 0.261188 0.0511875 0.336 ;
  RECT 0.0511875 0.240187 0.195562 0.261188 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.221812 0.066872 0.459375 0.0853125 ;
  RECT 0.221812 0.418687 0.459375 0.437063 ;
  RECT 0.459375 0.066872 0.494812 0.0853125 ;
  RECT 0.459375 0.418687 0.494812 0.437063 ;
  RECT 0.494812 0.066872 0.51319 0.0853125 ;
  RECT 0.494812 0.0853125 0.51319 0.418687 ;
  RECT 0.494812 0.418687 0.51319 0.437063 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.459375 0.522375 ;
  RECT 0.459375 0.485625 0.59456 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.59456 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.064969 0.0643125 0.0748125 0.122062 ;
  RECT 0.064969 0.122062 0.0748125 0.140437 ;
  RECT 0.0748125 0.0643125 0.093122 0.122062 ;
  RECT 0.0748125 0.122062 0.093122 0.140437 ;
  RECT 0.0748125 0.345845 0.093122 0.382595 ;
  RECT 0.0748125 0.382595 0.093122 0.439688 ;
  RECT 0.093122 0.0643125 0.103031 0.122062 ;
  RECT 0.093122 0.122062 0.103031 0.140437 ;
  RECT 0.093122 0.345845 0.103031 0.382595 ;
  RECT 0.103031 0.122062 0.232312 0.140437 ;
  RECT 0.103031 0.345845 0.232312 0.382595 ;
  RECT 0.232312 0.122062 0.250688 0.140437 ;
  RECT 0.232312 0.140437 0.250688 0.223781 ;
  RECT 0.232312 0.223781 0.250688 0.242156 ;
  RECT 0.232312 0.242156 0.250688 0.345845 ;
  RECT 0.232312 0.345845 0.250688 0.382595 ;
  RECT 0.250688 0.223781 0.459375 0.242156 ;
      LAYER M1 ;
  RECT 0.064969 0.0643125 0.0748125 0.122062 ;
  RECT 0.064969 0.122062 0.0748125 0.140437 ;
  RECT 0.0748125 0.0643125 0.093122 0.122062 ;
  RECT 0.0748125 0.122062 0.093122 0.140437 ;
  RECT 0.0748125 0.345845 0.093122 0.382595 ;
  RECT 0.0748125 0.382595 0.093122 0.439688 ;
  RECT 0.093122 0.0643125 0.103031 0.122062 ;
  RECT 0.093122 0.122062 0.103031 0.140437 ;
  RECT 0.093122 0.345845 0.103031 0.382595 ;
  RECT 0.103031 0.122062 0.232312 0.140437 ;
  RECT 0.103031 0.345845 0.232312 0.382595 ;
  RECT 0.232312 0.122062 0.250688 0.140437 ;
  RECT 0.232312 0.140437 0.250688 0.223781 ;
  RECT 0.232312 0.223781 0.250688 0.242156 ;
  RECT 0.232312 0.242156 0.250688 0.345845 ;
  RECT 0.232312 0.345845 0.250688 0.382595 ;
  RECT 0.250688 0.223781 0.459375 0.242156 ;
  END
END BUF_X8

MACRO BUF_X12
  CLASS core ;
  FOREIGN BUF_X12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.84 BY 0.504 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0315 0.154875 0.0525 0.240187 ;
  RECT 0.0315 0.240187 0.0525 0.261188 ;
  RECT 0.0315 0.261188 0.0525 0.33797 ;
  RECT 0.0525 0.240187 0.279562 0.261188 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.305812 0.066872 0.702185 0.0853125 ;
  RECT 0.305812 0.418687 0.702185 0.437063 ;
  RECT 0.702185 0.066872 0.745435 0.0853125 ;
  RECT 0.702185 0.418687 0.745435 0.437063 ;
  RECT 0.745435 0.066872 0.7665 0.0853125 ;
  RECT 0.745435 0.0853125 0.7665 0.418687 ;
  RECT 0.745435 0.418687 0.7665 0.437063 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.702185 0.522375 ;
  RECT 0.702185 0.485625 0.84656 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.84656 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0643125 0.361595 0.0735 0.382595 ;
  RECT 0.0643125 0.382595 0.0735 0.439688 ;
  RECT 0.0735 0.0643125 0.0945 0.121406 ;
  RECT 0.0735 0.121406 0.0945 0.142406 ;
  RECT 0.0735 0.361595 0.0945 0.382595 ;
  RECT 0.0735 0.382595 0.0945 0.439688 ;
  RECT 0.0945 0.121406 0.103031 0.142406 ;
  RECT 0.0945 0.361595 0.103031 0.382595 ;
  RECT 0.0945 0.382595 0.103031 0.439688 ;
  RECT 0.103031 0.121406 0.303187 0.142406 ;
  RECT 0.103031 0.361595 0.303187 0.382595 ;
  RECT 0.303187 0.121406 0.321562 0.142406 ;
  RECT 0.303187 0.142406 0.321562 0.242812 ;
  RECT 0.303187 0.242812 0.321562 0.261188 ;
  RECT 0.303187 0.261188 0.321562 0.361595 ;
  RECT 0.303187 0.361595 0.321562 0.382595 ;
  RECT 0.321562 0.242812 0.702185 0.261188 ;
      LAYER M1 ;
  RECT 0.0643125 0.361595 0.0735 0.382595 ;
  RECT 0.0643125 0.382595 0.0735 0.439688 ;
  RECT 0.0735 0.0643125 0.0945 0.121406 ;
  RECT 0.0735 0.121406 0.0945 0.142406 ;
  RECT 0.0735 0.361595 0.0945 0.382595 ;
  RECT 0.0735 0.382595 0.0945 0.439688 ;
  RECT 0.0945 0.121406 0.103031 0.142406 ;
  RECT 0.0945 0.361595 0.103031 0.382595 ;
  RECT 0.0945 0.382595 0.103031 0.439688 ;
  RECT 0.103031 0.121406 0.303187 0.142406 ;
  RECT 0.103031 0.361595 0.303187 0.382595 ;
  RECT 0.303187 0.121406 0.321562 0.142406 ;
  RECT 0.303187 0.142406 0.321562 0.242812 ;
  RECT 0.303187 0.242812 0.321562 0.261188 ;
  RECT 0.303187 0.261188 0.321562 0.361595 ;
  RECT 0.303187 0.361595 0.321562 0.382595 ;
  RECT 0.321562 0.242812 0.702185 0.261188 ;
  END
END BUF_X12

MACRO BUF_X16
  CLASS core ;
  FOREIGN BUF_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 1.092 BY 0.504 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.15225 0.0511875 0.232969 ;
  RECT 0.0328125 0.232969 0.0511875 0.27103 ;
  RECT 0.0328125 0.27103 0.0511875 0.336 ;
  RECT 0.0511875 0.232969 0.363563 0.27103 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.389813 0.066872 0.954185 0.0853125 ;
  RECT 0.389813 0.41475 0.954185 0.433125 ;
  RECT 0.954185 0.066872 0.9975 0.0853125 ;
  RECT 0.954185 0.41475 0.9975 0.433125 ;
  RECT 0.9975 0.066872 1.0185 0.0853125 ;
  RECT 0.9975 0.0853125 1.0185 0.41475 ;
  RECT 0.9975 0.41475 1.0185 0.433125 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.954185 0.522375 ;
  RECT 0.954185 0.485625 1.09856 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 1.09856 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0748125 0.0643125 0.093122 0.134531 ;
  RECT 0.0748125 0.134531 0.093122 0.152906 ;
  RECT 0.0748125 0.300563 0.093122 0.318937 ;
  RECT 0.0748125 0.318937 0.093122 0.42197 ;
  RECT 0.093122 0.134531 0.387188 0.152906 ;
  RECT 0.093122 0.300563 0.387188 0.318937 ;
  RECT 0.387188 0.134531 0.405562 0.152906 ;
  RECT 0.387188 0.152906 0.405562 0.2415 ;
  RECT 0.387188 0.2415 0.405562 0.259875 ;
  RECT 0.387188 0.259875 0.405562 0.300563 ;
  RECT 0.387188 0.300563 0.405562 0.318937 ;
  RECT 0.405562 0.2415 0.954185 0.259875 ;
      LAYER M1 ;
  RECT 0.0748125 0.0643125 0.093122 0.134531 ;
  RECT 0.0748125 0.134531 0.093122 0.152906 ;
  RECT 0.0748125 0.300563 0.093122 0.318937 ;
  RECT 0.0748125 0.318937 0.093122 0.42197 ;
  RECT 0.093122 0.134531 0.387188 0.152906 ;
  RECT 0.093122 0.300563 0.387188 0.318937 ;
  RECT 0.387188 0.134531 0.405562 0.152906 ;
  RECT 0.387188 0.152906 0.405562 0.2415 ;
  RECT 0.387188 0.2415 0.405562 0.259875 ;
  RECT 0.387188 0.259875 0.405562 0.300563 ;
  RECT 0.387188 0.300563 0.405562 0.318937 ;
  RECT 0.405562 0.2415 0.954185 0.259875 ;
  END
END BUF_X16

MACRO CLKBUF_X1
  CLASS core ;
  FOREIGN CLKBUF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.21 BY 0.504 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.126 0.0511875 0.378 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.1575 0.0748125 0.1785 0.462 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.093778 0.522375 ;
  RECT 0.093778 0.485625 0.216562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.216562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0748125 0.04725 0.075469 0.121406 ;
  RECT 0.0748125 0.121406 0.075469 0.139781 ;
  RECT 0.0748125 0.257905 0.075469 0.300563 ;
  RECT 0.0748125 0.300563 0.075469 0.34322 ;
  RECT 0.075469 0.04725 0.093122 0.121406 ;
  RECT 0.075469 0.121406 0.093122 0.139781 ;
  RECT 0.075469 0.139781 0.093122 0.257905 ;
  RECT 0.075469 0.257905 0.093122 0.300563 ;
  RECT 0.075469 0.300563 0.093122 0.34322 ;
  RECT 0.093122 0.121406 0.093778 0.139781 ;
  RECT 0.093122 0.139781 0.093778 0.257905 ;
  RECT 0.093122 0.257905 0.093778 0.300563 ;
      LAYER M1 ;
  RECT 0.0748125 0.04725 0.075469 0.121406 ;
  RECT 0.0748125 0.121406 0.075469 0.139781 ;
  RECT 0.0748125 0.257905 0.075469 0.300563 ;
  RECT 0.0748125 0.300563 0.075469 0.34322 ;
  RECT 0.075469 0.04725 0.093122 0.121406 ;
  RECT 0.075469 0.121406 0.093122 0.139781 ;
  RECT 0.075469 0.139781 0.093122 0.257905 ;
  RECT 0.075469 0.257905 0.093122 0.300563 ;
  RECT 0.075469 0.300563 0.093122 0.34322 ;
  RECT 0.093122 0.121406 0.093778 0.139781 ;
  RECT 0.093122 0.139781 0.093778 0.257905 ;
  RECT 0.093122 0.257905 0.093778 0.300563 ;
  END
END CLKBUF_X1

MACRO CLKBUF_X2
  CLASS core ;
  FOREIGN CLKBUF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.21 BY 0.504 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.19425 0.0511875 0.336 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.114122 0.418687 0.116812 0.462 ;
  RECT 0.116812 0.04725 0.135187 0.418687 ;
  RECT 0.116812 0.418687 0.135187 0.462 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.093122 0.522375 ;
  RECT 0.093122 0.485625 0.216562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.216562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0315 0.0846565 0.0525 0.126 ;
  RECT 0.0315 0.126 0.0525 0.144375 ;
  RECT 0.0315 0.364875 0.0525 0.38325 ;
  RECT 0.0315 0.38325 0.0525 0.450188 ;
  RECT 0.0525 0.126 0.0748125 0.144375 ;
  RECT 0.0525 0.364875 0.0748125 0.38325 ;
  RECT 0.0748125 0.126 0.093122 0.144375 ;
  RECT 0.0748125 0.144375 0.093122 0.364875 ;
  RECT 0.0748125 0.364875 0.093122 0.38325 ;
      LAYER M1 ;
  RECT 0.0315 0.0846565 0.0525 0.126 ;
  RECT 0.0315 0.126 0.0525 0.144375 ;
  RECT 0.0315 0.364875 0.0525 0.38325 ;
  RECT 0.0315 0.38325 0.0525 0.450188 ;
  RECT 0.0525 0.126 0.0748125 0.144375 ;
  RECT 0.0525 0.364875 0.0748125 0.38325 ;
  RECT 0.0748125 0.126 0.093122 0.144375 ;
  RECT 0.0748125 0.144375 0.093122 0.364875 ;
  RECT 0.0748125 0.364875 0.093122 0.38325 ;
  END
END CLKBUF_X2

MACRO CLKBUF_X4
  CLASS core ;
  FOREIGN CLKBUF_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.336 BY 0.504 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.158812 0.093122 0.345187 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.095156 0.066872 0.134531 0.0853125 ;
  RECT 0.134531 0.066872 0.135187 0.0853125 ;
  RECT 0.134531 0.418687 0.135187 0.437063 ;
  RECT 0.135187 0.066872 0.2415 0.0853125 ;
  RECT 0.135187 0.418687 0.2415 0.437063 ;
  RECT 0.2415 0.066872 0.2625 0.0853125 ;
  RECT 0.2415 0.0853125 0.2625 0.418687 ;
  RECT 0.2415 0.418687 0.2625 0.437063 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.135187 0.522375 ;
  RECT 0.135187 0.485625 0.342562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.342562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0269062 0.108937 0.0538125 0.127312 ;
  RECT 0.0538125 0.108937 0.116812 0.127312 ;
  RECT 0.0538125 0.376688 0.116812 0.395062 ;
  RECT 0.116812 0.108937 0.135187 0.127312 ;
  RECT 0.116812 0.127312 0.135187 0.376688 ;
  RECT 0.116812 0.376688 0.135187 0.395062 ;
      LAYER M1 ;
  RECT 0.0269062 0.108937 0.0538125 0.127312 ;
  RECT 0.0538125 0.108937 0.116812 0.127312 ;
  RECT 0.0538125 0.376688 0.116812 0.395062 ;
  RECT 0.116812 0.108937 0.135187 0.127312 ;
  RECT 0.116812 0.127312 0.135187 0.376688 ;
  RECT 0.116812 0.376688 0.135187 0.395062 ;
  END
END CLKBUF_X4

MACRO CLKBUF_X8
  CLASS core ;
  FOREIGN CLKBUF_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.588 BY 0.504 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.168 0.0511875 0.21525 ;
  RECT 0.0328125 0.21525 0.0511875 0.233625 ;
  RECT 0.0328125 0.233625 0.0511875 0.336 ;
  RECT 0.0511875 0.168 0.051844 0.21525 ;
  RECT 0.0511875 0.21525 0.051844 0.233625 ;
  RECT 0.051844 0.21525 0.208687 0.233625 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.221812 0.066872 0.471187 0.0853125 ;
  RECT 0.221812 0.418687 0.471187 0.437063 ;
  RECT 0.471187 0.066872 0.494812 0.0853125 ;
  RECT 0.471187 0.418687 0.494812 0.437063 ;
  RECT 0.494812 0.066872 0.51319 0.0853125 ;
  RECT 0.494812 0.0853125 0.51319 0.418687 ;
  RECT 0.494812 0.418687 0.51319 0.437063 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.471187 0.522375 ;
  RECT 0.471187 0.485625 0.59456 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.59456 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0328125 0.108937 0.0748125 0.127312 ;
  RECT 0.0748125 0.108937 0.093122 0.127312 ;
  RECT 0.0748125 0.295312 0.093122 0.316312 ;
  RECT 0.0748125 0.316312 0.093122 0.355687 ;
  RECT 0.093122 0.108937 0.266437 0.127312 ;
  RECT 0.093122 0.295312 0.266437 0.316312 ;
  RECT 0.266437 0.108937 0.284813 0.127312 ;
  RECT 0.266437 0.127312 0.284813 0.234281 ;
  RECT 0.266437 0.234281 0.284813 0.272345 ;
  RECT 0.266437 0.272345 0.284813 0.295312 ;
  RECT 0.266437 0.295312 0.284813 0.316312 ;
  RECT 0.284813 0.234281 0.471187 0.272345 ;
      LAYER M1 ;
  RECT 0.0328125 0.108937 0.0748125 0.127312 ;
  RECT 0.0748125 0.108937 0.093122 0.127312 ;
  RECT 0.0748125 0.295312 0.093122 0.316312 ;
  RECT 0.0748125 0.316312 0.093122 0.355687 ;
  RECT 0.093122 0.108937 0.266437 0.127312 ;
  RECT 0.093122 0.295312 0.266437 0.316312 ;
  RECT 0.266437 0.108937 0.284813 0.127312 ;
  RECT 0.266437 0.127312 0.284813 0.234281 ;
  RECT 0.266437 0.234281 0.284813 0.272345 ;
  RECT 0.266437 0.272345 0.284813 0.295312 ;
  RECT 0.266437 0.295312 0.284813 0.316312 ;
  RECT 0.284813 0.234281 0.471187 0.272345 ;
  END
END CLKBUF_X8

MACRO CLKBUF_X12
  CLASS core ;
  FOREIGN CLKBUF_X12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.84 BY 0.504 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0295312 0.156187 0.054469 0.2205 ;
  RECT 0.0295312 0.2205 0.054469 0.2415 ;
  RECT 0.0295312 0.2415 0.054469 0.347813 ;
  RECT 0.054469 0.2205 0.279562 0.2415 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.305812 0.066872 0.654935 0.0853125 ;
  RECT 0.305812 0.418687 0.654935 0.437063 ;
  RECT 0.654935 0.066872 0.745435 0.0853125 ;
  RECT 0.654935 0.418687 0.745435 0.437063 ;
  RECT 0.745435 0.066872 0.7665 0.0853125 ;
  RECT 0.745435 0.0853125 0.7665 0.418687 ;
  RECT 0.745435 0.418687 0.7665 0.437063 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.654935 0.522375 ;
  RECT 0.654935 0.485625 0.84656 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.84656 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.028153 0.108937 0.0748125 0.127312 ;
  RECT 0.0748125 0.108937 0.093122 0.127312 ;
  RECT 0.0748125 0.360938 0.093122 0.379312 ;
  RECT 0.0748125 0.379312 0.093122 0.439688 ;
  RECT 0.093122 0.108937 0.303187 0.127312 ;
  RECT 0.093122 0.360938 0.303187 0.379312 ;
  RECT 0.303187 0.108937 0.321562 0.127312 ;
  RECT 0.303187 0.127312 0.321562 0.206062 ;
  RECT 0.303187 0.206062 0.321562 0.226997 ;
  RECT 0.303187 0.226997 0.321562 0.360938 ;
  RECT 0.303187 0.360938 0.321562 0.379312 ;
  RECT 0.321562 0.108937 0.324188 0.127312 ;
  RECT 0.321562 0.127312 0.324188 0.206062 ;
  RECT 0.321562 0.206062 0.324188 0.226997 ;
  RECT 0.324188 0.206062 0.654935 0.226997 ;
      LAYER M1 ;
  RECT 0.028153 0.108937 0.0748125 0.127312 ;
  RECT 0.0748125 0.108937 0.093122 0.127312 ;
  RECT 0.0748125 0.360938 0.093122 0.379312 ;
  RECT 0.0748125 0.379312 0.093122 0.439688 ;
  RECT 0.093122 0.108937 0.303187 0.127312 ;
  RECT 0.093122 0.360938 0.303187 0.379312 ;
  RECT 0.303187 0.108937 0.321562 0.127312 ;
  RECT 0.303187 0.127312 0.321562 0.206062 ;
  RECT 0.303187 0.206062 0.321562 0.226997 ;
  RECT 0.303187 0.226997 0.321562 0.360938 ;
  RECT 0.303187 0.360938 0.321562 0.379312 ;
  RECT 0.321562 0.108937 0.324188 0.127312 ;
  RECT 0.321562 0.127312 0.324188 0.206062 ;
  RECT 0.321562 0.206062 0.324188 0.226997 ;
  RECT 0.324188 0.206062 0.654935 0.226997 ;
  END
END CLKBUF_X12

MACRO CLKBUF_X16
  CLASS core ;
  FOREIGN CLKBUF_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 1.092 BY 0.504 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.145687 0.0511875 0.213937 ;
  RECT 0.0328125 0.213937 0.0511875 0.234937 ;
  RECT 0.0328125 0.234937 0.0511875 0.345187 ;
  RECT 0.0511875 0.213937 0.363563 0.234937 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.389813 0.057028 0.954185 0.095156 ;
  RECT 0.389813 0.408845 0.954185 0.446905 ;
  RECT 0.954185 0.057028 0.9975 0.095156 ;
  RECT 0.954185 0.408845 0.9975 0.446905 ;
  RECT 0.9975 0.057028 1.0185 0.095156 ;
  RECT 0.9975 0.095156 1.0185 0.408845 ;
  RECT 0.9975 0.408845 1.0185 0.446905 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.954185 0.522375 ;
  RECT 0.954185 0.485625 1.09856 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 1.09856 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0748125 0.0715315 0.093122 0.134531 ;
  RECT 0.0748125 0.134531 0.093122 0.152906 ;
  RECT 0.0748125 0.34453 0.093122 0.369403 ;
  RECT 0.0748125 0.369403 0.093122 0.418687 ;
  RECT 0.093122 0.134531 0.39047 0.152906 ;
  RECT 0.093122 0.34453 0.39047 0.369403 ;
  RECT 0.39047 0.134531 0.42853 0.152906 ;
  RECT 0.39047 0.152906 0.42853 0.207375 ;
  RECT 0.39047 0.207375 0.42853 0.225684 ;
  RECT 0.39047 0.225684 0.42853 0.34453 ;
  RECT 0.39047 0.34453 0.42853 0.369403 ;
  RECT 0.42853 0.207375 0.954185 0.225684 ;
      LAYER M1 ;
  RECT 0.0748125 0.0715315 0.093122 0.134531 ;
  RECT 0.0748125 0.134531 0.093122 0.152906 ;
  RECT 0.0748125 0.34453 0.093122 0.369403 ;
  RECT 0.0748125 0.369403 0.093122 0.418687 ;
  RECT 0.093122 0.134531 0.39047 0.152906 ;
  RECT 0.093122 0.34453 0.39047 0.369403 ;
  RECT 0.39047 0.134531 0.42853 0.152906 ;
  RECT 0.39047 0.152906 0.42853 0.207375 ;
  RECT 0.39047 0.207375 0.42853 0.225684 ;
  RECT 0.39047 0.225684 0.42853 0.34453 ;
  RECT 0.39047 0.34453 0.42853 0.369403 ;
  RECT 0.42853 0.207375 0.954185 0.225684 ;
  END
END CLKBUF_X16

MACRO CLKGATETST_X1
  CLASS core ;
  FOREIGN CLKGATETST_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.714 BY 0.504 ;
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
  RECT 0.452748 0.156187 0.471187 0.336 ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.168 0.093122 0.441 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.21 0.0511875 0.441 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.662815 0.063 0.681185 0.429187 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.240187 0.522375 ;
  RECT 0.240187 0.485625 0.597185 0.522375 ;
  RECT 0.597185 0.485625 0.63919 0.522375 ;
  RECT 0.63919 0.485625 0.72056 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.72056 0.018375 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
  RECT 0.137812 0.263813 0.450188 0.282187 ;
  RECT 0.0958125 0.305812 0.342562 0.324188 ;
  RECT 0.479063 0.263813 0.66019 0.282187 ;
      LAYER MINT1 ;
  RECT 0.137812 0.263813 0.450188 0.282187 ;
  RECT 0.0958125 0.305812 0.342562 0.324188 ;
  RECT 0.479063 0.263813 0.66019 0.282187 ;
      LAYER M1 ;
  RECT 0.0315 0.066872 0.0525 0.0853125 ;
  RECT 0.0315 0.0853125 0.0525 0.139781 ;
  RECT 0.0525 0.066872 0.156187 0.0853125 ;
  RECT 0.158812 0.17325 0.177187 0.35503 ;
  RECT 0.242812 0.158812 0.261188 0.329437 ;
  RECT 0.303187 0.244125 0.324188 0.334688 ;
  RECT 0.410813 0.108937 0.429187 0.127312 ;
  RECT 0.410813 0.127312 0.429187 0.364875 ;
  RECT 0.410813 0.364875 0.429187 0.3885 ;
  RECT 0.429187 0.108937 0.492188 0.127312 ;
  RECT 0.429187 0.364875 0.492188 0.3885 ;
  RECT 0.492188 0.108937 0.49547 0.127312 ;
  RECT 0.494812 0.16275 0.518435 0.303845 ;
  RECT 0.494812 0.303845 0.518435 0.329437 ;
  RECT 0.518435 0.303845 0.53675 0.329437 ;
  RECT 0.53675 0.303845 0.555185 0.329437 ;
  RECT 0.53675 0.329437 0.555185 0.38325 ;
  RECT 0.62081 0.148312 0.63919 0.376688 ;
  RECT 0.116812 0.108937 0.135187 0.127312 ;
  RECT 0.116812 0.127312 0.135187 0.412125 ;
  RECT 0.116812 0.412125 0.135187 0.443625 ;
  RECT 0.135187 0.108937 0.198187 0.127312 ;
  RECT 0.135187 0.412125 0.198187 0.443625 ;
  RECT 0.198187 0.412125 0.240187 0.443625 ;
  RECT 0.200812 0.201469 0.219187 0.358312 ;
  RECT 0.200812 0.358312 0.219187 0.376688 ;
  RECT 0.219187 0.358312 0.366187 0.376688 ;
  RECT 0.366187 0.12075 0.387188 0.201469 ;
  RECT 0.366187 0.201469 0.387188 0.358312 ;
  RECT 0.366187 0.358312 0.387188 0.376688 ;
  RECT 0.284813 0.066872 0.303187 0.0853125 ;
  RECT 0.284813 0.0853125 0.303187 0.219187 ;
  RECT 0.303187 0.066872 0.305812 0.0853125 ;
  RECT 0.305812 0.066872 0.57881 0.0853125 ;
  RECT 0.305812 0.412125 0.57881 0.443625 ;
  RECT 0.57881 0.066872 0.597185 0.0853125 ;
  RECT 0.57881 0.0853125 0.597185 0.219187 ;
  RECT 0.57881 0.219187 0.597185 0.412125 ;
  RECT 0.57881 0.412125 0.597185 0.443625 ;
      LAYER V1 ;
  RECT 0.116812 0.305812 0.135187 0.324188 ;
  RECT 0.158812 0.263813 0.177187 0.282187 ;
  RECT 0.242812 0.263813 0.261188 0.282187 ;
  RECT 0.303187 0.305812 0.321562 0.324188 ;
  RECT 0.410813 0.263813 0.429187 0.282187 ;
  RECT 0.50006 0.263813 0.518435 0.282187 ;
  RECT 0.62081 0.263813 0.63919 0.282187 ;
      LAYER M1 ;
  RECT 0.0315 0.066872 0.0525 0.0853125 ;
  RECT 0.0315 0.0853125 0.0525 0.139781 ;
  RECT 0.0525 0.066872 0.156187 0.0853125 ;
  RECT 0.158812 0.17325 0.177187 0.35503 ;
  RECT 0.242812 0.158812 0.261188 0.329437 ;
  RECT 0.303187 0.244125 0.324188 0.334688 ;
  RECT 0.410813 0.108937 0.429187 0.127312 ;
  RECT 0.410813 0.127312 0.429187 0.364875 ;
  RECT 0.410813 0.364875 0.429187 0.3885 ;
  RECT 0.429187 0.108937 0.492188 0.127312 ;
  RECT 0.429187 0.364875 0.492188 0.3885 ;
  RECT 0.492188 0.108937 0.49547 0.127312 ;
  RECT 0.494812 0.16275 0.518435 0.303845 ;
  RECT 0.494812 0.303845 0.518435 0.329437 ;
  RECT 0.518435 0.303845 0.53675 0.329437 ;
  RECT 0.53675 0.303845 0.555185 0.329437 ;
  RECT 0.53675 0.329437 0.555185 0.38325 ;
  RECT 0.62081 0.148312 0.63919 0.376688 ;
  RECT 0.116812 0.108937 0.135187 0.127312 ;
  RECT 0.116812 0.127312 0.135187 0.412125 ;
  RECT 0.116812 0.412125 0.135187 0.443625 ;
  RECT 0.135187 0.108937 0.198187 0.127312 ;
  RECT 0.135187 0.412125 0.198187 0.443625 ;
  RECT 0.198187 0.412125 0.240187 0.443625 ;
  RECT 0.200812 0.201469 0.219187 0.358312 ;
  RECT 0.200812 0.358312 0.219187 0.376688 ;
  RECT 0.219187 0.358312 0.366187 0.376688 ;
  RECT 0.366187 0.12075 0.387188 0.201469 ;
  RECT 0.366187 0.201469 0.387188 0.358312 ;
  RECT 0.366187 0.358312 0.387188 0.376688 ;
  RECT 0.284813 0.066872 0.303187 0.0853125 ;
  RECT 0.284813 0.0853125 0.303187 0.219187 ;
  RECT 0.303187 0.066872 0.305812 0.0853125 ;
  RECT 0.305812 0.066872 0.57881 0.0853125 ;
  RECT 0.305812 0.412125 0.57881 0.443625 ;
  RECT 0.57881 0.066872 0.597185 0.0853125 ;
  RECT 0.57881 0.0853125 0.597185 0.219187 ;
  RECT 0.57881 0.219187 0.597185 0.412125 ;
  RECT 0.57881 0.412125 0.597185 0.443625 ;
  END
END CLKGATETST_X1

MACRO DFFRNQ_X1
  CLASS core ;
  FOREIGN DFFRNQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 1.092 BY 0.504 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.158812 0.177187 0.345187 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
  RECT 0.462 0.179812 0.744125 0.198187 ;
  RECT 0.744125 0.179812 0.87019 0.198187 ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.168 0.0511875 0.336 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 1.0395 0.042 1.0605 0.462 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.093122 0.522375 ;
  RECT 0.093122 0.485625 0.135187 0.522375 ;
  RECT 0.135187 0.485625 0.219187 0.522375 ;
  RECT 0.219187 0.485625 0.261188 0.522375 ;
  RECT 0.261188 0.485625 0.345187 0.522375 ;
  RECT 0.345187 0.485625 0.53412 0.522375 ;
  RECT 0.53412 0.485625 0.597185 0.522375 ;
  RECT 0.597185 0.485625 0.63919 0.522375 ;
  RECT 0.63919 0.485625 0.723185 0.522375 ;
  RECT 0.723185 0.485625 0.779625 0.522375 ;
  RECT 0.779625 0.485625 0.9765 0.522375 ;
  RECT 0.9765 0.485625 1.09856 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 1.09856 0.018375 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
  RECT 0.0958125 0.137812 0.744125 0.156187 ;
  RECT 0.0538125 0.347813 0.744125 0.366187 ;
      LAYER MINT1 ;
  RECT 0.0958125 0.137812 0.744125 0.156187 ;
  RECT 0.0538125 0.347813 0.744125 0.366187 ;
      LAYER M1 ;
  RECT 0.116812 0.04725 0.135187 0.456685 ;
  RECT 0.200812 0.04725 0.219187 0.456685 ;
  RECT 0.347813 0.408845 0.53412 0.446905 ;
  RECT 0.284813 0.066872 0.303187 0.0853125 ;
  RECT 0.284813 0.0853125 0.303187 0.287438 ;
  RECT 0.284813 0.287438 0.303187 0.439688 ;
  RECT 0.303187 0.066872 0.525 0.0853125 ;
  RECT 0.525 0.066872 0.543375 0.0853125 ;
  RECT 0.525 0.0853125 0.543375 0.287438 ;
  RECT 0.378 0.216562 0.396375 0.332062 ;
  RECT 0.378 0.332062 0.396375 0.350438 ;
  RECT 0.396375 0.332062 0.57881 0.350438 ;
  RECT 0.57881 0.04725 0.597185 0.216562 ;
  RECT 0.57881 0.216562 0.597185 0.332062 ;
  RECT 0.57881 0.332062 0.597185 0.350438 ;
  RECT 0.57881 0.350438 0.597185 0.441 ;
  RECT 0.662815 0.066872 0.681185 0.0853125 ;
  RECT 0.662815 0.0853125 0.681185 0.240187 ;
  RECT 0.662815 0.240187 0.681185 0.439688 ;
  RECT 0.681185 0.066872 0.876095 0.0853125 ;
  RECT 0.876095 0.066872 0.89447 0.0853125 ;
  RECT 0.876095 0.0853125 0.89447 0.240187 ;
  RECT 0.80325 0.258562 0.821625 0.418687 ;
  RECT 0.80325 0.418687 0.821625 0.437063 ;
  RECT 0.821625 0.418687 0.95681 0.437063 ;
  RECT 0.95681 0.04725 0.975185 0.086625 ;
  RECT 0.95681 0.086625 0.975185 0.258562 ;
  RECT 0.95681 0.258562 0.975185 0.418687 ;
  RECT 0.95681 0.418687 0.975185 0.437063 ;
  RECT 0.975185 0.086625 0.9765 0.258562 ;
  RECT 0.975185 0.258562 0.9765 0.418687 ;
  RECT 0.975185 0.418687 0.9765 0.437063 ;
  RECT 0.0315 0.055781 0.0525 0.0924655 ;
  RECT 0.0315 0.0924655 0.0525 0.110906 ;
  RECT 0.0315 0.372028 0.0525 0.397688 ;
  RECT 0.0315 0.397688 0.0525 0.450188 ;
  RECT 0.0525 0.0924655 0.0748125 0.110906 ;
  RECT 0.0525 0.372028 0.0748125 0.397688 ;
  RECT 0.0748125 0.0924655 0.093122 0.110906 ;
  RECT 0.0748125 0.110906 0.093122 0.372028 ;
  RECT 0.0748125 0.372028 0.093122 0.397688 ;
  RECT 0.242812 0.127312 0.261188 0.324188 ;
  RECT 0.326813 0.263813 0.345187 0.376688 ;
  RECT 0.345187 0.127312 0.366187 0.192937 ;
  RECT 0.483 0.169312 0.501375 0.287438 ;
  RECT 0.62081 0.179812 0.63919 0.379312 ;
  RECT 0.70481 0.114122 0.723185 0.208031 ;
  RECT 0.70481 0.301875 0.723185 0.408187 ;
  RECT 0.758625 0.108937 0.779625 0.450188 ;
  RECT 0.83081 0.114122 0.849185 0.208687 ;
      LAYER V1 ;
  RECT 0.0748125 0.347813 0.093122 0.366187 ;
  RECT 0.116812 0.137812 0.135187 0.156187 ;
  RECT 0.242812 0.137812 0.261188 0.156187 ;
  RECT 0.326813 0.347813 0.345187 0.366187 ;
  RECT 0.347813 0.137812 0.366187 0.156187 ;
  RECT 0.483 0.179812 0.501375 0.198187 ;
  RECT 0.62081 0.347813 0.63919 0.366187 ;
  RECT 0.70481 0.137812 0.723185 0.156187 ;
  RECT 0.70481 0.347813 0.723185 0.366187 ;
  RECT 0.83081 0.179812 0.849185 0.198187 ;
      LAYER M1 ;
  RECT 0.116812 0.04725 0.135187 0.456685 ;
  RECT 0.200812 0.04725 0.219187 0.456685 ;
  RECT 0.347813 0.408845 0.53412 0.446905 ;
  RECT 0.284813 0.066872 0.303187 0.0853125 ;
  RECT 0.284813 0.0853125 0.303187 0.287438 ;
  RECT 0.284813 0.287438 0.303187 0.439688 ;
  RECT 0.303187 0.066872 0.525 0.0853125 ;
  RECT 0.525 0.066872 0.543375 0.0853125 ;
  RECT 0.525 0.0853125 0.543375 0.287438 ;
  RECT 0.378 0.216562 0.396375 0.332062 ;
  RECT 0.378 0.332062 0.396375 0.350438 ;
  RECT 0.396375 0.332062 0.57881 0.350438 ;
  RECT 0.57881 0.04725 0.597185 0.216562 ;
  RECT 0.57881 0.216562 0.597185 0.332062 ;
  RECT 0.57881 0.332062 0.597185 0.350438 ;
  RECT 0.57881 0.350438 0.597185 0.441 ;
  RECT 0.662815 0.066872 0.681185 0.0853125 ;
  RECT 0.662815 0.0853125 0.681185 0.240187 ;
  RECT 0.662815 0.240187 0.681185 0.439688 ;
  RECT 0.681185 0.066872 0.876095 0.0853125 ;
  RECT 0.876095 0.066872 0.89447 0.0853125 ;
  RECT 0.876095 0.0853125 0.89447 0.240187 ;
  RECT 0.80325 0.258562 0.821625 0.418687 ;
  RECT 0.80325 0.418687 0.821625 0.437063 ;
  RECT 0.821625 0.418687 0.95681 0.437063 ;
  RECT 0.95681 0.04725 0.975185 0.086625 ;
  RECT 0.95681 0.086625 0.975185 0.258562 ;
  RECT 0.95681 0.258562 0.975185 0.418687 ;
  RECT 0.95681 0.418687 0.975185 0.437063 ;
  RECT 0.975185 0.086625 0.9765 0.258562 ;
  RECT 0.975185 0.258562 0.9765 0.418687 ;
  RECT 0.975185 0.418687 0.9765 0.437063 ;
  RECT 0.0315 0.055781 0.0525 0.0924655 ;
  RECT 0.0315 0.0924655 0.0525 0.110906 ;
  RECT 0.0315 0.372028 0.0525 0.397688 ;
  RECT 0.0315 0.397688 0.0525 0.450188 ;
  RECT 0.0525 0.0924655 0.0748125 0.110906 ;
  RECT 0.0525 0.372028 0.0748125 0.397688 ;
  RECT 0.0748125 0.0924655 0.093122 0.110906 ;
  RECT 0.0748125 0.110906 0.093122 0.372028 ;
  RECT 0.0748125 0.372028 0.093122 0.397688 ;
  RECT 0.242812 0.127312 0.261188 0.324188 ;
  RECT 0.326813 0.263813 0.345187 0.376688 ;
  RECT 0.345187 0.127312 0.366187 0.192937 ;
  RECT 0.483 0.169312 0.501375 0.287438 ;
  RECT 0.62081 0.179812 0.63919 0.379312 ;
  RECT 0.70481 0.114122 0.723185 0.208031 ;
  RECT 0.70481 0.301875 0.723185 0.408187 ;
  RECT 0.758625 0.108937 0.779625 0.450188 ;
  RECT 0.83081 0.114122 0.849185 0.208687 ;
  END
END DFFRNQ_X1

MACRO DFFSNQ_X1
  CLASS core ;
  FOREIGN DFFSNQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 1.092 BY 0.504 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.158812 0.177187 0.345187 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
  RECT 0.473813 0.179812 0.744125 0.198187 ;
  RECT 0.744125 0.179812 0.87019 0.198187 ;
    END
  END SN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.168 0.0511875 0.336 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 1.0395 0.042 1.0605 0.462 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.093122 0.522375 ;
  RECT 0.093122 0.485625 0.135187 0.522375 ;
  RECT 0.135187 0.485625 0.219187 0.522375 ;
  RECT 0.219187 0.485625 0.261188 0.522375 ;
  RECT 0.261188 0.485625 0.345187 0.522375 ;
  RECT 0.345187 0.485625 0.363563 0.522375 ;
  RECT 0.363563 0.485625 0.597185 0.522375 ;
  RECT 0.597185 0.485625 0.63919 0.522375 ;
  RECT 0.63919 0.485625 0.72581 0.522375 ;
  RECT 0.72581 0.485625 0.91212 0.522375 ;
  RECT 0.91212 0.485625 0.9765 0.522375 ;
  RECT 0.9765 0.485625 1.09856 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 1.09856 0.018375 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
  RECT 0.0958125 0.137812 0.744125 0.156187 ;
  RECT 0.0538125 0.347813 0.744125 0.366187 ;
      LAYER MINT1 ;
  RECT 0.0958125 0.137812 0.744125 0.156187 ;
  RECT 0.0538125 0.347813 0.744125 0.366187 ;
      LAYER M1 ;
  RECT 0.116812 0.04725 0.135187 0.456685 ;
  RECT 0.200812 0.04725 0.219187 0.456685 ;
  RECT 0.284813 0.0800625 0.303187 0.0984375 ;
  RECT 0.284813 0.0984375 0.303187 0.240187 ;
  RECT 0.284813 0.240187 0.303187 0.439688 ;
  RECT 0.303187 0.0800625 0.53675 0.0984375 ;
  RECT 0.53675 0.0800625 0.555185 0.0984375 ;
  RECT 0.53675 0.0984375 0.555185 0.240187 ;
  RECT 0.62081 0.179812 0.63919 0.376688 ;
  RECT 0.70481 0.127312 0.72581 0.213281 ;
  RECT 0.70481 0.257905 0.72581 0.389813 ;
  RECT 0.83081 0.122062 0.849185 0.208687 ;
  RECT 0.788815 0.258562 0.807185 0.376688 ;
  RECT 0.788815 0.376688 0.807185 0.395062 ;
  RECT 0.807185 0.376688 0.95681 0.395062 ;
  RECT 0.95681 0.04725 0.975185 0.086625 ;
  RECT 0.95681 0.086625 0.975185 0.258562 ;
  RECT 0.95681 0.258562 0.975185 0.376688 ;
  RECT 0.95681 0.376688 0.975185 0.395062 ;
  RECT 0.975185 0.086625 0.9765 0.258562 ;
  RECT 0.975185 0.258562 0.9765 0.376688 ;
  RECT 0.975185 0.376688 0.9765 0.395062 ;
  RECT 0.0295312 0.0538125 0.0315 0.0905625 ;
  RECT 0.0295312 0.0905625 0.0315 0.116156 ;
  RECT 0.0315 0.0538125 0.0525 0.0905625 ;
  RECT 0.0315 0.0905625 0.0525 0.116156 ;
  RECT 0.0315 0.372028 0.0525 0.397688 ;
  RECT 0.0315 0.397688 0.0525 0.450188 ;
  RECT 0.0525 0.0538125 0.054469 0.0905625 ;
  RECT 0.0525 0.0905625 0.054469 0.116156 ;
  RECT 0.0525 0.372028 0.054469 0.397688 ;
  RECT 0.054469 0.0905625 0.0748125 0.116156 ;
  RECT 0.054469 0.372028 0.0748125 0.397688 ;
  RECT 0.0748125 0.0905625 0.093122 0.116156 ;
  RECT 0.0748125 0.116156 0.093122 0.372028 ;
  RECT 0.0748125 0.372028 0.093122 0.397688 ;
  RECT 0.242812 0.127312 0.261188 0.324188 ;
  RECT 0.326813 0.263813 0.345187 0.387188 ;
  RECT 0.345187 0.127312 0.363563 0.200156 ;
  RECT 0.494812 0.169312 0.51319 0.240187 ;
  RECT 0.399 0.179812 0.417375 0.376688 ;
  RECT 0.399 0.376688 0.417375 0.395062 ;
  RECT 0.417375 0.376688 0.576185 0.395062 ;
  RECT 0.576185 0.376688 0.57881 0.395062 ;
  RECT 0.576185 0.395062 0.57881 0.450188 ;
  RECT 0.57881 0.063 0.597185 0.179812 ;
  RECT 0.57881 0.179812 0.597185 0.376688 ;
  RECT 0.57881 0.376688 0.597185 0.395062 ;
  RECT 0.57881 0.395062 0.597185 0.450188 ;
  RECT 0.662815 0.0748125 0.681185 0.093122 ;
  RECT 0.662815 0.093122 0.681185 0.240187 ;
  RECT 0.662815 0.240187 0.681185 0.441 ;
  RECT 0.681185 0.0748125 0.88725 0.093122 ;
  RECT 0.88725 0.0748125 0.90556 0.093122 ;
  RECT 0.88725 0.093122 0.90556 0.240187 ;
  RECT 0.72581 0.418687 0.91212 0.437063 ;
      LAYER V1 ;
  RECT 0.0748125 0.347813 0.093122 0.366187 ;
  RECT 0.116812 0.137812 0.135187 0.156187 ;
  RECT 0.242812 0.137812 0.261188 0.156187 ;
  RECT 0.326813 0.347813 0.345187 0.366187 ;
  RECT 0.345187 0.137812 0.363563 0.156187 ;
  RECT 0.494812 0.179812 0.51319 0.198187 ;
  RECT 0.62081 0.347813 0.63919 0.366187 ;
  RECT 0.70481 0.137812 0.723185 0.156187 ;
  RECT 0.70481 0.347813 0.723185 0.366187 ;
  RECT 0.83081 0.179812 0.849185 0.198187 ;
      LAYER M1 ;
  RECT 0.116812 0.04725 0.135187 0.456685 ;
  RECT 0.200812 0.04725 0.219187 0.456685 ;
  RECT 0.284813 0.0800625 0.303187 0.0984375 ;
  RECT 0.284813 0.0984375 0.303187 0.240187 ;
  RECT 0.284813 0.240187 0.303187 0.439688 ;
  RECT 0.303187 0.0800625 0.53675 0.0984375 ;
  RECT 0.53675 0.0800625 0.555185 0.0984375 ;
  RECT 0.53675 0.0984375 0.555185 0.240187 ;
  RECT 0.62081 0.179812 0.63919 0.376688 ;
  RECT 0.70481 0.127312 0.72581 0.213281 ;
  RECT 0.70481 0.257905 0.72581 0.389813 ;
  RECT 0.83081 0.122062 0.849185 0.208687 ;
  RECT 0.788815 0.258562 0.807185 0.376688 ;
  RECT 0.788815 0.376688 0.807185 0.395062 ;
  RECT 0.807185 0.376688 0.95681 0.395062 ;
  RECT 0.95681 0.04725 0.975185 0.086625 ;
  RECT 0.95681 0.086625 0.975185 0.258562 ;
  RECT 0.95681 0.258562 0.975185 0.376688 ;
  RECT 0.95681 0.376688 0.975185 0.395062 ;
  RECT 0.975185 0.086625 0.9765 0.258562 ;
  RECT 0.975185 0.258562 0.9765 0.376688 ;
  RECT 0.975185 0.376688 0.9765 0.395062 ;
  RECT 0.0295312 0.0538125 0.0315 0.0905625 ;
  RECT 0.0295312 0.0905625 0.0315 0.116156 ;
  RECT 0.0315 0.0538125 0.0525 0.0905625 ;
  RECT 0.0315 0.0905625 0.0525 0.116156 ;
  RECT 0.0315 0.372028 0.0525 0.397688 ;
  RECT 0.0315 0.397688 0.0525 0.450188 ;
  RECT 0.0525 0.0538125 0.054469 0.0905625 ;
  RECT 0.0525 0.0905625 0.054469 0.116156 ;
  RECT 0.0525 0.372028 0.054469 0.397688 ;
  RECT 0.054469 0.0905625 0.0748125 0.116156 ;
  RECT 0.054469 0.372028 0.0748125 0.397688 ;
  RECT 0.0748125 0.0905625 0.093122 0.116156 ;
  RECT 0.0748125 0.116156 0.093122 0.372028 ;
  RECT 0.0748125 0.372028 0.093122 0.397688 ;
  RECT 0.242812 0.127312 0.261188 0.324188 ;
  RECT 0.326813 0.263813 0.345187 0.387188 ;
  RECT 0.345187 0.127312 0.363563 0.200156 ;
  RECT 0.494812 0.169312 0.51319 0.240187 ;
  RECT 0.399 0.179812 0.417375 0.376688 ;
  RECT 0.399 0.376688 0.417375 0.395062 ;
  RECT 0.417375 0.376688 0.576185 0.395062 ;
  RECT 0.576185 0.376688 0.57881 0.395062 ;
  RECT 0.576185 0.395062 0.57881 0.450188 ;
  RECT 0.57881 0.063 0.597185 0.179812 ;
  RECT 0.57881 0.179812 0.597185 0.376688 ;
  RECT 0.57881 0.376688 0.597185 0.395062 ;
  RECT 0.57881 0.395062 0.597185 0.450188 ;
  RECT 0.662815 0.0748125 0.681185 0.093122 ;
  RECT 0.662815 0.093122 0.681185 0.240187 ;
  RECT 0.662815 0.240187 0.681185 0.441 ;
  RECT 0.681185 0.0748125 0.88725 0.093122 ;
  RECT 0.88725 0.0748125 0.90556 0.093122 ;
  RECT 0.88725 0.093122 0.90556 0.240187 ;
  RECT 0.72581 0.418687 0.91212 0.437063 ;
  END
END DFFSNQ_X1

MACRO FA_X1
  CLASS core ;
  FOREIGN FA_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 1.008 BY 0.504 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
  RECT 0.137812 0.305812 0.72056 0.324188 ;
      LAYER V1 ;
  RECT 0.4305 0.305812 0.448875 0.324188 ;
  RECT 0.681185 0.305812 0.69956 0.324188 ;
      LAYER M1 ;
  RECT 0.4305 0.263813 0.448875 0.345187 ;
  RECT 0.681185 0.179812 0.70481 0.345187 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
  RECT 0.179812 0.179812 0.51778 0.198187 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
  RECT 0.0958125 0.137812 0.828185 0.156187 ;
      LAYER V1 ;
  RECT 0.116812 0.137812 0.135187 0.156187 ;
  RECT 0.380625 0.137812 0.399 0.156187 ;
  RECT 0.788815 0.137812 0.807185 0.156187 ;
      LAYER M1 ;
  RECT 0.116812 0.127312 0.135187 0.387188 ;
  RECT 0.380625 0.127312 0.399 0.240187 ;
  RECT 0.788815 0.116812 0.807185 0.240187 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.95681 0.0748125 0.975185 0.429187 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.53675 0.135844 0.555185 0.42 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.093122 0.522375 ;
  RECT 0.093122 0.485625 0.177187 0.522375 ;
  RECT 0.177187 0.485625 0.219187 0.522375 ;
  RECT 0.219187 0.485625 0.4305 0.522375 ;
  RECT 0.4305 0.485625 0.503345 0.522375 ;
  RECT 0.503345 0.485625 0.681185 0.522375 ;
  RECT 0.681185 0.485625 0.711375 0.522375 ;
  RECT 0.711375 0.485625 0.76519 0.522375 ;
  RECT 0.76519 0.485625 0.845905 0.522375 ;
  RECT 0.845905 0.485625 0.89119 0.522375 ;
  RECT 0.89119 0.485625 1.01456 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 1.01456 0.018375 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
  RECT 0.0538125 0.263813 0.866905 0.282187 ;
  RECT 0.263813 0.221812 0.91212 0.240187 ;
      LAYER MINT1 ;
  RECT 0.0538125 0.263813 0.866905 0.282187 ;
  RECT 0.263813 0.221812 0.91212 0.240187 ;
      LAYER M1 ;
  RECT 0.0177187 0.116812 0.0426562 0.221812 ;
  RECT 0.0177187 0.221812 0.0426562 0.240187 ;
  RECT 0.0426562 0.221812 0.0675935 0.240187 ;
  RECT 0.0675935 0.221812 0.093122 0.240187 ;
  RECT 0.0675935 0.240187 0.093122 0.303187 ;
  RECT 0.158812 0.179812 0.177187 0.387188 ;
  RECT 0.27825 0.179812 0.303187 0.33272 ;
  RECT 0.242812 0.063656 0.405562 0.0885935 ;
  RECT 0.242812 0.377345 0.263813 0.39572 ;
  RECT 0.242812 0.39572 0.263813 0.457998 ;
  RECT 0.263813 0.377345 0.4095 0.39572 ;
  RECT 0.4095 0.377345 0.4305 0.39572 ;
  RECT 0.4095 0.39572 0.4305 0.457998 ;
  RECT 0.4095 0.457998 0.4305 0.462 ;
  RECT 0.478405 0.160125 0.503345 0.3045 ;
  RECT 0.57881 0.127312 0.597185 0.240187 ;
  RECT 0.57881 0.368812 0.597185 0.387188 ;
  RECT 0.57881 0.387188 0.597185 0.456685 ;
  RECT 0.597185 0.368812 0.662815 0.387188 ;
  RECT 0.662815 0.368812 0.681185 0.387188 ;
  RECT 0.662815 0.387188 0.681185 0.456685 ;
  RECT 0.74675 0.04725 0.76519 0.456685 ;
  RECT 0.827465 0.253312 0.845905 0.387188 ;
  RECT 0.200812 0.063 0.219187 0.441 ;
  RECT 0.326813 0.179812 0.345187 0.33272 ;
  RECT 0.62081 0.179812 0.64575 0.324188 ;
  RECT 0.555185 0.065625 0.711375 0.086625 ;
  RECT 0.87281 0.179812 0.89119 0.345187 ;
      LAYER V1 ;
  RECT 0.0748125 0.263813 0.093122 0.282187 ;
  RECT 0.158812 0.305812 0.177187 0.324188 ;
  RECT 0.200812 0.179812 0.219187 0.198187 ;
  RECT 0.284813 0.221812 0.303187 0.240187 ;
  RECT 0.326813 0.263813 0.345187 0.282187 ;
  RECT 0.478405 0.179812 0.49678 0.198187 ;
  RECT 0.57881 0.137812 0.597185 0.156187 ;
  RECT 0.627375 0.263813 0.64575 0.282187 ;
  RECT 0.74675 0.221812 0.76519 0.240187 ;
  RECT 0.827465 0.263813 0.845905 0.282187 ;
  RECT 0.87281 0.221812 0.89119 0.240187 ;
      LAYER M1 ;
  RECT 0.0177187 0.116812 0.0426562 0.221812 ;
  RECT 0.0177187 0.221812 0.0426562 0.240187 ;
  RECT 0.0426562 0.221812 0.0675935 0.240187 ;
  RECT 0.0675935 0.221812 0.093122 0.240187 ;
  RECT 0.0675935 0.240187 0.093122 0.303187 ;
  RECT 0.158812 0.179812 0.177187 0.387188 ;
  RECT 0.27825 0.179812 0.303187 0.33272 ;
  RECT 0.242812 0.063656 0.405562 0.0885935 ;
  RECT 0.242812 0.377345 0.263813 0.39572 ;
  RECT 0.242812 0.39572 0.263813 0.457998 ;
  RECT 0.263813 0.377345 0.4095 0.39572 ;
  RECT 0.4095 0.377345 0.4305 0.39572 ;
  RECT 0.4095 0.39572 0.4305 0.457998 ;
  RECT 0.4095 0.457998 0.4305 0.462 ;
  RECT 0.478405 0.160125 0.503345 0.3045 ;
  RECT 0.57881 0.127312 0.597185 0.240187 ;
  RECT 0.57881 0.368812 0.597185 0.387188 ;
  RECT 0.57881 0.387188 0.597185 0.456685 ;
  RECT 0.597185 0.368812 0.662815 0.387188 ;
  RECT 0.662815 0.368812 0.681185 0.387188 ;
  RECT 0.662815 0.387188 0.681185 0.456685 ;
  RECT 0.74675 0.04725 0.76519 0.456685 ;
  RECT 0.827465 0.253312 0.845905 0.387188 ;
  RECT 0.200812 0.063 0.219187 0.441 ;
  RECT 0.326813 0.179812 0.345187 0.33272 ;
  RECT 0.62081 0.179812 0.64575 0.324188 ;
  RECT 0.555185 0.065625 0.711375 0.086625 ;
  RECT 0.87281 0.179812 0.89119 0.345187 ;
  END
END FA_X1

MACRO FILLTIE
  CLASS core ;
  FOREIGN FILLTIE 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.379312 BY 0.504 ;
  OBS
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.385875 0.018375 ;
  RECT -0.0065625 0.485625 0.385875 0.522375 ;
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.385875 0.018375 ;
  RECT -0.0065625 0.485625 0.385875 0.522375 ;
  END
END FILLTIE

MACRO FILL_X1
  CLASS core ;
  FOREIGN FILL_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.084 BY 0.504 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.0905625 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.0905625 0.018375 ;
    END
  END VSS
END FILL_X1

MACRO FILL_X2
  CLASS core ;
  FOREIGN FILL_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.126 BY 0.504 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.132562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.132562 0.018375 ;
    END
  END VSS
END FILL_X2

MACRO FILL_X4
  CLASS core ;
  FOREIGN FILL_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.21 BY 0.504 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.216562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.216562 0.018375 ;
    END
  END VSS
END FILL_X4

MACRO FILL_X8
  CLASS core ;
  FOREIGN FILL_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.378 BY 0.504 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.384562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.384562 0.018375 ;
    END
  END VSS
END FILL_X8

MACRO FILL_X16
  CLASS core ;
  FOREIGN FILL_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.714 BY 0.504 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.72056 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.72056 0.018375 ;
    END
  END VSS
END FILL_X16

MACRO HA_X1
  CLASS core ;
  FOREIGN HA_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.546 BY 0.504 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.179812 0.177187 0.364875 ;
  RECT 0.158812 0.364875 0.177187 0.38325 ;
  RECT 0.177187 0.364875 0.284813 0.38325 ;
  RECT 0.284813 0.179812 0.303187 0.364875 ;
  RECT 0.284813 0.364875 0.303187 0.38325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.200812 0.168 0.219187 0.336 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.0538125 0.0511875 0.418687 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.494812 0.118125 0.51319 0.418687 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.391125 0.522375 ;
  RECT 0.391125 0.485625 0.433125 0.522375 ;
  RECT 0.433125 0.485625 0.55256 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.55256 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.221812 0.066872 0.408187 0.0853125 ;
  RECT 0.266437 0.12075 0.326813 0.14175 ;
  RECT 0.326813 0.12075 0.347813 0.14175 ;
  RECT 0.326813 0.14175 0.347813 0.303187 ;
  RECT 0.326813 0.303187 0.347813 0.395062 ;
  RECT 0.347813 0.12075 0.41475 0.14175 ;
  RECT 0.41475 0.12075 0.433125 0.14175 ;
  RECT 0.41475 0.14175 0.433125 0.303187 ;
  RECT 0.0748125 0.108937 0.093122 0.129937 ;
  RECT 0.0748125 0.129937 0.093122 0.179812 ;
  RECT 0.0748125 0.179812 0.093122 0.418687 ;
  RECT 0.0748125 0.418687 0.093122 0.437063 ;
  RECT 0.093122 0.108937 0.242812 0.129937 ;
  RECT 0.093122 0.418687 0.242812 0.437063 ;
  RECT 0.242812 0.418687 0.371372 0.437063 ;
  RECT 0.371372 0.179812 0.391125 0.418687 ;
  RECT 0.371372 0.418687 0.391125 0.437063 ;
      LAYER M1 ;
  RECT 0.221812 0.066872 0.408187 0.0853125 ;
  RECT 0.266437 0.12075 0.326813 0.14175 ;
  RECT 0.326813 0.12075 0.347813 0.14175 ;
  RECT 0.326813 0.14175 0.347813 0.303187 ;
  RECT 0.326813 0.303187 0.347813 0.395062 ;
  RECT 0.347813 0.12075 0.41475 0.14175 ;
  RECT 0.41475 0.12075 0.433125 0.14175 ;
  RECT 0.41475 0.14175 0.433125 0.303187 ;
  RECT 0.0748125 0.108937 0.093122 0.129937 ;
  RECT 0.0748125 0.129937 0.093122 0.179812 ;
  RECT 0.0748125 0.179812 0.093122 0.418687 ;
  RECT 0.0748125 0.418687 0.093122 0.437063 ;
  RECT 0.093122 0.108937 0.242812 0.129937 ;
  RECT 0.093122 0.418687 0.242812 0.437063 ;
  RECT 0.242812 0.418687 0.371372 0.437063 ;
  RECT 0.371372 0.179812 0.391125 0.418687 ;
  RECT 0.371372 0.418687 0.391125 0.437063 ;
  END
END HA_X1

MACRO INV_X1
  CLASS core ;
  FOREIGN INV_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.126 BY 0.504 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.126 0.0511875 0.378 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.0748125 0.093122 0.42 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.132562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.132562 0.018375 ;
    END
  END VSS
END INV_X1

MACRO INV_X2
  CLASS core ;
  FOREIGN INV_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.168 BY 0.504 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.126 0.0511875 0.378 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.0853125 0.093122 0.378 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.174562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.174562 0.018375 ;
    END
  END VSS
END INV_X2

MACRO INV_X4
  CLASS core ;
  FOREIGN INV_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.504 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0315 0.168 0.0525 0.2415 ;
  RECT 0.0315 0.2415 0.0525 0.259875 ;
  RECT 0.0315 0.259875 0.0525 0.336 ;
  RECT 0.0525 0.2415 0.156187 0.259875 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0269062 0.093122 0.0387188 0.13125 ;
  RECT 0.0387188 0.093122 0.200812 0.13125 ;
  RECT 0.0387188 0.372685 0.200812 0.410813 ;
  RECT 0.200812 0.093122 0.219187 0.13125 ;
  RECT 0.200812 0.13125 0.219187 0.372685 ;
  RECT 0.200812 0.372685 0.219187 0.410813 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.258562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.258562 0.018375 ;
    END
  END VSS
END INV_X4

MACRO INV_X8
  CLASS core ;
  FOREIGN INV_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.42 BY 0.504 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.127312 0.093122 0.259875 ;
  RECT 0.0748125 0.259875 0.093122 0.298595 ;
  RECT 0.0748125 0.298595 0.093122 0.378 ;
  RECT 0.093122 0.259875 0.303187 0.298595 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0269062 0.414095 0.0354375 0.43247 ;
  RECT 0.0354375 0.0721875 0.36553 0.0905625 ;
  RECT 0.0354375 0.414095 0.36553 0.43247 ;
  RECT 0.36553 0.0721875 0.39047 0.0905625 ;
  RECT 0.36553 0.0905625 0.39047 0.414095 ;
  RECT 0.36553 0.414095 0.39047 0.43247 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.426563 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.426563 0.018375 ;
    END
  END VSS
END INV_X8

MACRO INV_X12
  CLASS core ;
  FOREIGN INV_X12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.588 BY 0.504 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.126 0.093122 0.2415 ;
  RECT 0.0748125 0.2415 0.093122 0.259875 ;
  RECT 0.0748125 0.259875 0.093122 0.378 ;
  RECT 0.093122 0.2415 0.450188 0.259875 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0354375 0.066872 0.533465 0.0853125 ;
  RECT 0.0354375 0.417375 0.533465 0.438375 ;
  RECT 0.533465 0.066872 0.55847 0.0853125 ;
  RECT 0.533465 0.0853125 0.55847 0.417375 ;
  RECT 0.533465 0.417375 0.55847 0.438375 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.59456 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.59456 0.018375 ;
    END
  END VSS
END INV_X12

MACRO INV_X16
  CLASS core ;
  FOREIGN INV_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.756 BY 0.504 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.168 0.0511875 0.242812 ;
  RECT 0.0328125 0.242812 0.0511875 0.261188 ;
  RECT 0.0328125 0.261188 0.0511875 0.369403 ;
  RECT 0.0511875 0.242812 0.61819 0.261188 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.702185 0.522375 ;
  RECT 0.702185 0.485625 0.762565 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.762565 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0354375 0.065625 0.681185 0.086625 ;
  RECT 0.0354375 0.408187 0.681185 0.446905 ;
  RECT 0.681185 0.065625 0.702185 0.086625 ;
  RECT 0.681185 0.086625 0.702185 0.408187 ;
  RECT 0.681185 0.408187 0.702185 0.446905 ;
      LAYER M1 ;
  RECT 0.0354375 0.065625 0.681185 0.086625 ;
  RECT 0.0354375 0.408187 0.681185 0.446905 ;
  RECT 0.681185 0.065625 0.702185 0.086625 ;
  RECT 0.681185 0.086625 0.702185 0.408187 ;
  RECT 0.681185 0.408187 0.702185 0.446905 ;
  END
END INV_X16

MACRO LHQ_X1
  CLASS core ;
  FOREIGN LHQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.588 BY 0.504 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.105 0.177187 0.336 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.168 0.0511875 0.336 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.53675 0.0853125 0.555185 0.418687 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.51319 0.522375 ;
  RECT 0.51319 0.485625 0.59456 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.59456 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0315 0.364875 0.0328125 0.38325 ;
  RECT 0.0315 0.38325 0.0328125 0.462 ;
  RECT 0.0328125 0.042 0.0511875 0.060375 ;
  RECT 0.0328125 0.060375 0.0511875 0.12075 ;
  RECT 0.0328125 0.12075 0.0511875 0.139125 ;
  RECT 0.0328125 0.364875 0.0511875 0.38325 ;
  RECT 0.0328125 0.38325 0.0511875 0.462 ;
  RECT 0.0511875 0.042 0.0525 0.060375 ;
  RECT 0.0511875 0.12075 0.0525 0.139125 ;
  RECT 0.0511875 0.364875 0.0525 0.38325 ;
  RECT 0.0511875 0.38325 0.0525 0.462 ;
  RECT 0.0525 0.042 0.0748125 0.060375 ;
  RECT 0.0525 0.12075 0.0748125 0.139125 ;
  RECT 0.0525 0.364875 0.0748125 0.38325 ;
  RECT 0.0748125 0.042 0.093122 0.060375 ;
  RECT 0.0748125 0.12075 0.093122 0.139125 ;
  RECT 0.0748125 0.139125 0.093122 0.211312 ;
  RECT 0.0748125 0.211312 0.093122 0.229687 ;
  RECT 0.0748125 0.229687 0.093122 0.271688 ;
  RECT 0.0748125 0.271688 0.093122 0.364875 ;
  RECT 0.0748125 0.364875 0.093122 0.38325 ;
  RECT 0.093122 0.042 0.212625 0.060375 ;
  RECT 0.212625 0.042 0.231 0.060375 ;
  RECT 0.212625 0.060375 0.231 0.12075 ;
  RECT 0.212625 0.12075 0.231 0.139125 ;
  RECT 0.212625 0.139125 0.231 0.211312 ;
  RECT 0.212625 0.211312 0.231 0.229687 ;
  RECT 0.231 0.211312 0.242812 0.229687 ;
  RECT 0.242812 0.211312 0.261188 0.229687 ;
  RECT 0.242812 0.229687 0.261188 0.271688 ;
  RECT 0.347813 0.0748125 0.366187 0.093122 ;
  RECT 0.347813 0.093122 0.366187 0.324188 ;
  RECT 0.366187 0.0748125 0.452748 0.093122 ;
  RECT 0.452748 0.0748125 0.471187 0.093122 ;
  RECT 0.452748 0.093122 0.471187 0.324188 ;
  RECT 0.452748 0.324188 0.471187 0.389155 ;
  RECT 0.116812 0.08925 0.135187 0.301875 ;
  RECT 0.116812 0.301875 0.135187 0.364875 ;
  RECT 0.116812 0.364875 0.135187 0.38325 ;
  RECT 0.135187 0.364875 0.200812 0.38325 ;
  RECT 0.200812 0.301875 0.223125 0.364875 ;
  RECT 0.200812 0.364875 0.223125 0.38325 ;
  RECT 0.179812 0.418687 0.254625 0.437063 ;
  RECT 0.254625 0.0748125 0.305812 0.113466 ;
  RECT 0.254625 0.418687 0.305812 0.437063 ;
  RECT 0.305812 0.0748125 0.324188 0.113466 ;
  RECT 0.305812 0.113466 0.324188 0.200812 ;
  RECT 0.305812 0.200812 0.324188 0.41803 ;
  RECT 0.305812 0.41803 0.324188 0.418687 ;
  RECT 0.305812 0.418687 0.324188 0.437063 ;
  RECT 0.324188 0.41803 0.494812 0.418687 ;
  RECT 0.324188 0.418687 0.494812 0.437063 ;
  RECT 0.494812 0.200812 0.51319 0.41803 ;
  RECT 0.494812 0.41803 0.51319 0.418687 ;
  RECT 0.494812 0.418687 0.51319 0.437063 ;
      LAYER M1 ;
  RECT 0.0315 0.364875 0.0328125 0.38325 ;
  RECT 0.0315 0.38325 0.0328125 0.462 ;
  RECT 0.0328125 0.042 0.0511875 0.060375 ;
  RECT 0.0328125 0.060375 0.0511875 0.12075 ;
  RECT 0.0328125 0.12075 0.0511875 0.139125 ;
  RECT 0.0328125 0.364875 0.0511875 0.38325 ;
  RECT 0.0328125 0.38325 0.0511875 0.462 ;
  RECT 0.0511875 0.042 0.0525 0.060375 ;
  RECT 0.0511875 0.12075 0.0525 0.139125 ;
  RECT 0.0511875 0.364875 0.0525 0.38325 ;
  RECT 0.0511875 0.38325 0.0525 0.462 ;
  RECT 0.0525 0.042 0.0748125 0.060375 ;
  RECT 0.0525 0.12075 0.0748125 0.139125 ;
  RECT 0.0525 0.364875 0.0748125 0.38325 ;
  RECT 0.0748125 0.042 0.093122 0.060375 ;
  RECT 0.0748125 0.12075 0.093122 0.139125 ;
  RECT 0.0748125 0.139125 0.093122 0.211312 ;
  RECT 0.0748125 0.211312 0.093122 0.229687 ;
  RECT 0.0748125 0.229687 0.093122 0.271688 ;
  RECT 0.0748125 0.271688 0.093122 0.364875 ;
  RECT 0.0748125 0.364875 0.093122 0.38325 ;
  RECT 0.093122 0.042 0.212625 0.060375 ;
  RECT 0.212625 0.042 0.231 0.060375 ;
  RECT 0.212625 0.060375 0.231 0.12075 ;
  RECT 0.212625 0.12075 0.231 0.139125 ;
  RECT 0.212625 0.139125 0.231 0.211312 ;
  RECT 0.212625 0.211312 0.231 0.229687 ;
  RECT 0.231 0.211312 0.242812 0.229687 ;
  RECT 0.242812 0.211312 0.261188 0.229687 ;
  RECT 0.242812 0.229687 0.261188 0.271688 ;
  RECT 0.347813 0.0748125 0.366187 0.093122 ;
  RECT 0.347813 0.093122 0.366187 0.324188 ;
  RECT 0.366187 0.0748125 0.452748 0.093122 ;
  RECT 0.452748 0.0748125 0.471187 0.093122 ;
  RECT 0.452748 0.093122 0.471187 0.324188 ;
  RECT 0.452748 0.324188 0.471187 0.389155 ;
  RECT 0.116812 0.08925 0.135187 0.301875 ;
  RECT 0.116812 0.301875 0.135187 0.364875 ;
  RECT 0.116812 0.364875 0.135187 0.38325 ;
  RECT 0.135187 0.364875 0.200812 0.38325 ;
  RECT 0.200812 0.301875 0.223125 0.364875 ;
  RECT 0.200812 0.364875 0.223125 0.38325 ;
  RECT 0.179812 0.418687 0.254625 0.437063 ;
  RECT 0.254625 0.0748125 0.305812 0.113466 ;
  RECT 0.254625 0.418687 0.305812 0.437063 ;
  RECT 0.305812 0.0748125 0.324188 0.113466 ;
  RECT 0.305812 0.113466 0.324188 0.200812 ;
  RECT 0.305812 0.200812 0.324188 0.41803 ;
  RECT 0.305812 0.41803 0.324188 0.418687 ;
  RECT 0.305812 0.418687 0.324188 0.437063 ;
  RECT 0.324188 0.41803 0.494812 0.418687 ;
  RECT 0.324188 0.418687 0.494812 0.437063 ;
  RECT 0.494812 0.200812 0.51319 0.41803 ;
  RECT 0.494812 0.41803 0.51319 0.418687 ;
  RECT 0.494812 0.418687 0.51319 0.437063 ;
  END
END LHQ_X1

MACRO MUX2_X1
  CLASS core ;
  FOREIGN MUX2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.546 BY 0.504 ;
  PIN I0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.368812 0.158812 0.387188 0.345187 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.168 0.093122 0.294 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
  RECT 0.0774375 0.431812 0.258562 0.450188 ;
      LAYER V1 ;
  RECT 0.0984375 0.431812 0.135187 0.450188 ;
      LAYER M1 ;
  RECT 0.0177187 0.158812 0.0360938 0.431812 ;
  RECT 0.0177187 0.431812 0.0360938 0.450188 ;
  RECT 0.0360938 0.431812 0.145687 0.450188 ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.452748 0.126 0.471187 0.418687 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.303187 0.522375 ;
  RECT 0.303187 0.485625 0.345187 0.522375 ;
  RECT 0.345187 0.485625 0.51319 0.522375 ;
  RECT 0.51319 0.485625 0.55256 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.55256 0.018375 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
  RECT 0.179812 0.221812 0.366187 0.240187 ;
      LAYER MINT1 ;
  RECT 0.179812 0.221812 0.366187 0.240187 ;
      LAYER M1 ;
  RECT 0.0525 0.106312 0.064969 0.124687 ;
  RECT 0.064969 0.106312 0.103031 0.124687 ;
  RECT 0.064969 0.322875 0.103031 0.34125 ;
  RECT 0.064969 0.34125 0.103031 0.378 ;
  RECT 0.103031 0.106312 0.200812 0.124687 ;
  RECT 0.103031 0.322875 0.200812 0.34125 ;
  RECT 0.200812 0.106312 0.219187 0.124687 ;
  RECT 0.200812 0.124687 0.219187 0.322875 ;
  RECT 0.200812 0.322875 0.219187 0.34125 ;
  RECT 0.190312 0.431812 0.284813 0.462 ;
  RECT 0.284813 0.200812 0.303187 0.431812 ;
  RECT 0.284813 0.431812 0.303187 0.462 ;
  RECT 0.326813 0.179812 0.345187 0.280875 ;
  RECT 0.242812 0.057028 0.261188 0.0958125 ;
  RECT 0.242812 0.0958125 0.261188 0.324188 ;
  RECT 0.242812 0.324188 0.261188 0.402938 ;
  RECT 0.261188 0.057028 0.494812 0.0958125 ;
  RECT 0.494812 0.057028 0.51319 0.0958125 ;
  RECT 0.494812 0.0958125 0.51319 0.324188 ;
      LAYER V1 ;
  RECT 0.200812 0.221812 0.219187 0.240187 ;
  RECT 0.200812 0.431812 0.237562 0.450188 ;
  RECT 0.326813 0.221812 0.345187 0.240187 ;
      LAYER M1 ;
  RECT 0.0525 0.106312 0.064969 0.124687 ;
  RECT 0.064969 0.106312 0.103031 0.124687 ;
  RECT 0.064969 0.322875 0.103031 0.34125 ;
  RECT 0.064969 0.34125 0.103031 0.378 ;
  RECT 0.103031 0.106312 0.200812 0.124687 ;
  RECT 0.103031 0.322875 0.200812 0.34125 ;
  RECT 0.200812 0.106312 0.219187 0.124687 ;
  RECT 0.200812 0.124687 0.219187 0.322875 ;
  RECT 0.200812 0.322875 0.219187 0.34125 ;
  RECT 0.190312 0.431812 0.284813 0.462 ;
  RECT 0.284813 0.200812 0.303187 0.431812 ;
  RECT 0.284813 0.431812 0.303187 0.462 ;
  RECT 0.326813 0.179812 0.345187 0.280875 ;
  RECT 0.242812 0.057028 0.261188 0.0958125 ;
  RECT 0.242812 0.0958125 0.261188 0.324188 ;
  RECT 0.242812 0.324188 0.261188 0.402938 ;
  RECT 0.261188 0.057028 0.494812 0.0958125 ;
  RECT 0.494812 0.057028 0.51319 0.0958125 ;
  RECT 0.494812 0.0958125 0.51319 0.324188 ;
  END
END MUX2_X1

MACRO NAND2_X1
  CLASS core ;
  FOREIGN NAND2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.168 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.168 0.135187 0.376688 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.168 0.0511875 0.376688 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.0872815 0.093122 0.126 ;
  RECT 0.0748125 0.126 0.093122 0.418687 ;
  RECT 0.093122 0.0872815 0.1155 0.126 ;
  RECT 0.1155 0.042 0.1365 0.0872815 ;
  RECT 0.1155 0.0872815 0.1365 0.126 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.174562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.174562 0.018375 ;
    END
  END VSS
END NAND2_X1

MACRO NAND2_X2
  CLASS core ;
  FOREIGN NAND2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.147656 0.135187 0.362905 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.179812 0.0511875 0.443625 ;
  RECT 0.0328125 0.443625 0.0511875 0.462 ;
  RECT 0.0511875 0.443625 0.200812 0.462 ;
  RECT 0.200812 0.179812 0.219187 0.443625 ;
  RECT 0.200812 0.443625 0.219187 0.462 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.080719 0.093122 0.118781 ;
  RECT 0.0748125 0.118781 0.093122 0.27825 ;
  RECT 0.0748125 0.27825 0.093122 0.39178 ;
  RECT 0.0748125 0.39178 0.093122 0.42 ;
  RECT 0.093122 0.080719 0.158812 0.118781 ;
  RECT 0.093122 0.39178 0.158812 0.42 ;
  RECT 0.158812 0.080719 0.177187 0.118781 ;
  RECT 0.158812 0.27825 0.177187 0.39178 ;
  RECT 0.158812 0.39178 0.177187 0.42 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.258562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.258562 0.018375 ;
    END
  END VSS
END NAND2_X2

MACRO NAND3_X1
  CLASS core ;
  FOREIGN NAND3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.21 0.177187 0.294 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.167344 0.135187 0.336 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.141094 0.0511875 0.376688 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.0538125 0.093122 0.0721875 ;
  RECT 0.0748125 0.0721875 0.093122 0.168 ;
  RECT 0.0748125 0.168 0.093122 0.336 ;
  RECT 0.0748125 0.336 0.093122 0.443625 ;
  RECT 0.0748125 0.443625 0.093122 0.462 ;
  RECT 0.093122 0.0538125 0.158812 0.0721875 ;
  RECT 0.093122 0.443625 0.158812 0.462 ;
  RECT 0.158812 0.042 0.1995 0.0538125 ;
  RECT 0.158812 0.0538125 0.1995 0.0721875 ;
  RECT 0.158812 0.443625 0.1995 0.462 ;
  RECT 0.1995 0.042 0.200812 0.0538125 ;
  RECT 0.1995 0.0538125 0.200812 0.0721875 ;
  RECT 0.1995 0.0721875 0.200812 0.168 ;
  RECT 0.1995 0.443625 0.200812 0.462 ;
  RECT 0.200812 0.042 0.219187 0.0538125 ;
  RECT 0.200812 0.0538125 0.219187 0.0721875 ;
  RECT 0.200812 0.0721875 0.219187 0.168 ;
  RECT 0.200812 0.336 0.219187 0.443625 ;
  RECT 0.200812 0.443625 0.219187 0.462 ;
  RECT 0.219187 0.042 0.2205 0.0538125 ;
  RECT 0.219187 0.0538125 0.2205 0.0721875 ;
  RECT 0.219187 0.0721875 0.2205 0.168 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.258562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.258562 0.018375 ;
    END
  END VSS
END NAND3_X1

MACRO NAND3_X2
  CLASS core ;
  FOREIGN NAND3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.378 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.326813 0.21 0.345187 0.336 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.197531 0.163406 0.222469 0.336 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.168 0.093122 0.336 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0177187 0.372685 0.240187 0.410813 ;
  RECT 0.240187 0.372685 0.284813 0.410813 ;
  RECT 0.284813 0.122062 0.303187 0.372685 ;
  RECT 0.284813 0.372685 0.303187 0.410813 ;
  RECT 0.303187 0.372685 0.324188 0.410813 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.240187 0.522375 ;
  RECT 0.240187 0.485625 0.345187 0.522375 ;
  RECT 0.345187 0.485625 0.384562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.384562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.137812 0.0728435 0.326813 0.0924655 ;
  RECT 0.326813 0.0728435 0.345187 0.0924655 ;
  RECT 0.326813 0.0924655 0.345187 0.147656 ;
  RECT 0.0328125 0.116156 0.240187 0.137156 ;
      LAYER M1 ;
  RECT 0.137812 0.0728435 0.326813 0.0924655 ;
  RECT 0.326813 0.0728435 0.345187 0.0924655 ;
  RECT 0.326813 0.0924655 0.345187 0.147656 ;
  RECT 0.0328125 0.116156 0.240187 0.137156 ;
  END
END NAND3_X2

MACRO NAND4_X1
  CLASS core ;
  FOREIGN NAND4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.242812 0.168 0.261188 0.376688 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.158812 0.177187 0.336 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.127312 0.135187 0.294 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.127312 0.0511875 0.376688 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.336 0.093122 0.42328 ;
  RECT 0.0748125 0.42328 0.093122 0.462 ;
  RECT 0.093122 0.42328 0.200812 0.462 ;
  RECT 0.200812 0.107625 0.219187 0.126 ;
  RECT 0.200812 0.126 0.219187 0.336 ;
  RECT 0.200812 0.336 0.219187 0.42328 ;
  RECT 0.200812 0.42328 0.219187 0.462 ;
  RECT 0.219187 0.107625 0.239531 0.126 ;
  RECT 0.239531 0.042 0.26447 0.107625 ;
  RECT 0.239531 0.107625 0.26447 0.126 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.300563 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.300563 0.018375 ;
    END
  END VSS
END NAND4_X1

MACRO NAND4_X2
  CLASS core ;
  FOREIGN NAND4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.462 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.366187 0.234937 0.389813 0.336 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.242812 0.223125 0.261188 0.345187 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.158812 0.135187 0.336 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.168656 0.0511875 0.336 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0735 0.36422 0.0945 0.378 ;
  RECT 0.0735 0.378 0.0945 0.418687 ;
  RECT 0.0735 0.418687 0.0945 0.437063 ;
  RECT 0.0945 0.418687 0.284813 0.437063 ;
  RECT 0.284813 0.192937 0.303187 0.211312 ;
  RECT 0.284813 0.211312 0.303187 0.359625 ;
  RECT 0.284813 0.359625 0.303187 0.36422 ;
  RECT 0.284813 0.36422 0.303187 0.378 ;
  RECT 0.284813 0.418687 0.303187 0.437063 ;
  RECT 0.303187 0.192937 0.368812 0.211312 ;
  RECT 0.303187 0.359625 0.368812 0.36422 ;
  RECT 0.303187 0.36422 0.368812 0.378 ;
  RECT 0.303187 0.418687 0.368812 0.437063 ;
  RECT 0.368812 0.192937 0.387188 0.211312 ;
  RECT 0.368812 0.359625 0.387188 0.36422 ;
  RECT 0.368812 0.36422 0.387188 0.378 ;
  RECT 0.368812 0.378 0.387188 0.418687 ;
  RECT 0.368812 0.418687 0.387188 0.437063 ;
  RECT 0.387188 0.192937 0.429187 0.211312 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.4305 0.522375 ;
  RECT 0.4305 0.485625 0.468562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.468562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0315 0.066872 0.0525 0.0853125 ;
  RECT 0.0315 0.0853125 0.0525 0.139781 ;
  RECT 0.0525 0.066872 0.282187 0.0853125 ;
  RECT 0.179812 0.150937 0.4095 0.169312 ;
  RECT 0.4095 0.042 0.4305 0.150937 ;
  RECT 0.4095 0.150937 0.4305 0.169312 ;
  RECT 0.0958125 0.108937 0.324188 0.127312 ;
      LAYER M1 ;
  RECT 0.0315 0.066872 0.0525 0.0853125 ;
  RECT 0.0315 0.0853125 0.0525 0.139781 ;
  RECT 0.0525 0.066872 0.282187 0.0853125 ;
  RECT 0.179812 0.150937 0.4095 0.169312 ;
  RECT 0.4095 0.042 0.4305 0.150937 ;
  RECT 0.4095 0.150937 0.4305 0.169312 ;
  RECT 0.0958125 0.108937 0.324188 0.127312 ;
  END
END NAND4_X2

MACRO NOR2_X1
  CLASS core ;
  FOREIGN NOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.168 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.127312 0.135187 0.336 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.127312 0.0511875 0.336 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.0853125 0.093122 0.378 ;
  RECT 0.0748125 0.378 0.093122 0.41672 ;
  RECT 0.093122 0.378 0.1155 0.41672 ;
  RECT 0.1155 0.378 0.1365 0.41672 ;
  RECT 0.1155 0.41672 0.1365 0.462 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.174562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.174562 0.018375 ;
    END
  END VSS
END NOR2_X1

MACRO NOR2_X2
  CLASS core ;
  FOREIGN NOR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.141094 0.135187 0.336 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.042 0.0511875 0.060375 ;
  RECT 0.0328125 0.060375 0.0511875 0.324188 ;
  RECT 0.0511875 0.042 0.200812 0.060375 ;
  RECT 0.200812 0.042 0.219187 0.060375 ;
  RECT 0.200812 0.060375 0.219187 0.324188 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.084 0.093122 0.102375 ;
  RECT 0.0748125 0.102375 0.093122 0.225684 ;
  RECT 0.0748125 0.225684 0.093122 0.364875 ;
  RECT 0.0748125 0.364875 0.093122 0.38325 ;
  RECT 0.093122 0.084 0.1155 0.102375 ;
  RECT 0.093122 0.364875 0.1155 0.38325 ;
  RECT 0.1155 0.084 0.1365 0.102375 ;
  RECT 0.1155 0.364875 0.1365 0.38325 ;
  RECT 0.1155 0.38325 0.1365 0.42 ;
  RECT 0.1365 0.084 0.158812 0.102375 ;
  RECT 0.158812 0.084 0.177187 0.102375 ;
  RECT 0.158812 0.102375 0.177187 0.225684 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.258562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.258562 0.018375 ;
    END
  END VSS
END NOR2_X2

MACRO NOR3_X1
  CLASS core ;
  FOREIGN NOR3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.21 0.177187 0.294 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.127312 0.135187 0.362905 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.127312 0.0511875 0.362905 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.042 0.093122 0.060375 ;
  RECT 0.0748125 0.060375 0.093122 0.168 ;
  RECT 0.0748125 0.168 0.093122 0.336 ;
  RECT 0.0748125 0.336 0.093122 0.402938 ;
  RECT 0.0748125 0.402938 0.093122 0.421312 ;
  RECT 0.093122 0.042 0.198844 0.060375 ;
  RECT 0.093122 0.402938 0.198844 0.421312 ;
  RECT 0.198844 0.042 0.1995 0.060375 ;
  RECT 0.198844 0.060375 0.1995 0.168 ;
  RECT 0.198844 0.402938 0.1995 0.421312 ;
  RECT 0.1995 0.042 0.2205 0.060375 ;
  RECT 0.1995 0.060375 0.2205 0.168 ;
  RECT 0.1995 0.336 0.2205 0.402938 ;
  RECT 0.1995 0.402938 0.2205 0.421312 ;
  RECT 0.1995 0.421312 0.2205 0.462 ;
  RECT 0.2205 0.042 0.221156 0.060375 ;
  RECT 0.2205 0.060375 0.221156 0.168 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.258562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.258562 0.018375 ;
    END
  END VSS
END NOR3_X1

MACRO NOR3_X2
  CLASS core ;
  FOREIGN NOR3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.378 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.326813 0.168 0.345187 0.294 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.200812 0.168 0.219187 0.336655 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.168 0.0511875 0.340595 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.056372 0.101062 0.284813 0.139125 ;
  RECT 0.284813 0.101062 0.303187 0.139125 ;
  RECT 0.284813 0.139125 0.303187 0.378 ;
  RECT 0.303187 0.101062 0.321562 0.139125 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.345187 0.522375 ;
  RECT 0.345187 0.485625 0.384562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.384562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.137812 0.41147 0.326813 0.429845 ;
  RECT 0.326813 0.338625 0.345187 0.41147 ;
  RECT 0.326813 0.41147 0.345187 0.429845 ;
  RECT 0.056372 0.36553 0.249375 0.387845 ;
      LAYER M1 ;
  RECT 0.137812 0.41147 0.326813 0.429845 ;
  RECT 0.326813 0.338625 0.345187 0.41147 ;
  RECT 0.326813 0.41147 0.345187 0.429845 ;
  RECT 0.056372 0.36553 0.249375 0.387845 ;
  END
END NOR3_X2

MACRO NOR4_X1
  CLASS core ;
  FOREIGN NOR4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.242812 0.127312 0.261188 0.336 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.127312 0.177187 0.336 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.168 0.135187 0.376688 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.127312 0.0511875 0.376688 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.042 0.093122 0.066872 ;
  RECT 0.0748125 0.066872 0.093122 0.141094 ;
  RECT 0.093122 0.042 0.200812 0.066872 ;
  RECT 0.200812 0.042 0.219187 0.066872 ;
  RECT 0.200812 0.066872 0.219187 0.141094 ;
  RECT 0.200812 0.141094 0.219187 0.378 ;
  RECT 0.200812 0.378 0.219187 0.396375 ;
  RECT 0.219187 0.378 0.239531 0.396375 ;
  RECT 0.239531 0.378 0.26447 0.396375 ;
  RECT 0.239531 0.396375 0.26447 0.462 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.300563 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.300563 0.018375 ;
    END
  END VSS
END NOR4_X1

MACRO NOR4_X2
  CLASS core ;
  FOREIGN NOR4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.462 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.366187 0.168 0.389813 0.266437 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.242812 0.158812 0.261188 0.287438 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.158812 0.177187 0.345187 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.168 0.135187 0.338625 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0735 0.066872 0.0945 0.0853125 ;
  RECT 0.0735 0.0853125 0.0945 0.126 ;
  RECT 0.0735 0.126 0.0945 0.139781 ;
  RECT 0.0945 0.066872 0.284813 0.0853125 ;
  RECT 0.284813 0.066872 0.303187 0.0853125 ;
  RECT 0.284813 0.126 0.303187 0.139781 ;
  RECT 0.284813 0.139781 0.303187 0.144375 ;
  RECT 0.284813 0.144375 0.303187 0.290063 ;
  RECT 0.284813 0.290063 0.303187 0.308437 ;
  RECT 0.303187 0.066872 0.368812 0.0853125 ;
  RECT 0.303187 0.126 0.368812 0.139781 ;
  RECT 0.303187 0.139781 0.368812 0.144375 ;
  RECT 0.303187 0.290063 0.368812 0.308437 ;
  RECT 0.368812 0.066872 0.387188 0.0853125 ;
  RECT 0.368812 0.0853125 0.387188 0.126 ;
  RECT 0.368812 0.126 0.387188 0.139781 ;
  RECT 0.368812 0.139781 0.387188 0.144375 ;
  RECT 0.368812 0.290063 0.387188 0.308437 ;
  RECT 0.387188 0.290063 0.435095 0.308437 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.282187 0.522375 ;
  RECT 0.282187 0.485625 0.324188 0.522375 ;
  RECT 0.324188 0.485625 0.4305 0.522375 ;
  RECT 0.4305 0.485625 0.468562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.468562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.137812 0.373997 0.324188 0.395062 ;
  RECT 0.0315 0.36422 0.0525 0.418687 ;
  RECT 0.0315 0.418687 0.0525 0.437063 ;
  RECT 0.0525 0.418687 0.282187 0.437063 ;
  RECT 0.221812 0.332062 0.4095 0.350438 ;
  RECT 0.4095 0.332062 0.4305 0.350438 ;
  RECT 0.4095 0.350438 0.4305 0.450188 ;
      LAYER M1 ;
  RECT 0.137812 0.373997 0.324188 0.395062 ;
  RECT 0.0315 0.36422 0.0525 0.418687 ;
  RECT 0.0315 0.418687 0.0525 0.437063 ;
  RECT 0.0525 0.418687 0.282187 0.437063 ;
  RECT 0.221812 0.332062 0.4095 0.350438 ;
  RECT 0.4095 0.332062 0.4305 0.350438 ;
  RECT 0.4095 0.350438 0.4305 0.450188 ;
  END
END NOR4_X2

MACRO OAI21_X1
  CLASS core ;
  FOREIGN OAI21_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.168 0.135187 0.378 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.168 0.0511875 0.416063 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.200812 0.168 0.219187 0.378 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.168 0.093122 0.417375 ;
  RECT 0.0748125 0.417375 0.093122 0.438375 ;
  RECT 0.093122 0.417375 0.195562 0.438375 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.195562 0.522375 ;
  RECT 0.195562 0.485625 0.258562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.258562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0328125 0.0479062 0.0511875 0.101719 ;
  RECT 0.0328125 0.101719 0.0511875 0.122719 ;
  RECT 0.0511875 0.101719 0.195562 0.122719 ;
      LAYER M1 ;
  RECT 0.0328125 0.0479062 0.0511875 0.101719 ;
  RECT 0.0328125 0.101719 0.0511875 0.122719 ;
  RECT 0.0511875 0.101719 0.195562 0.122719 ;
  END
END OAI21_X1

MACRO OAI21_X2
  CLASS core ;
  FOREIGN OAI21_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.378 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.239531 0.21 0.26447 0.294 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.158812 0.177187 0.185653 ;
  RECT 0.158812 0.185653 0.177187 0.329437 ;
  RECT 0.158812 0.329437 0.177187 0.347813 ;
  RECT 0.177187 0.329437 0.326813 0.347813 ;
  RECT 0.326813 0.185653 0.345187 0.329437 ;
  RECT 0.326813 0.329437 0.345187 0.347813 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.168 0.093122 0.34453 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0190312 0.373997 0.116812 0.395062 ;
  RECT 0.116812 0.108937 0.135187 0.127312 ;
  RECT 0.116812 0.127312 0.135187 0.182437 ;
  RECT 0.116812 0.182437 0.135187 0.373997 ;
  RECT 0.116812 0.373997 0.135187 0.395062 ;
  RECT 0.135187 0.108937 0.279562 0.127312 ;
  RECT 0.135187 0.373997 0.279562 0.395062 ;
  RECT 0.279562 0.108937 0.284813 0.127312 ;
  RECT 0.284813 0.108937 0.303187 0.127312 ;
  RECT 0.284813 0.127312 0.303187 0.182437 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.351095 0.522375 ;
  RECT 0.351095 0.485625 0.384562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.384562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0315 0.066872 0.0525 0.0853125 ;
  RECT 0.0315 0.0853125 0.0525 0.139781 ;
  RECT 0.0525 0.066872 0.326813 0.0853125 ;
  RECT 0.326813 0.066872 0.345187 0.0853125 ;
  RECT 0.326813 0.0853125 0.345187 0.139781 ;
  RECT 0.326813 0.139781 0.345187 0.141094 ;
  RECT 0.0958125 0.418687 0.351095 0.437063 ;
      LAYER M1 ;
  RECT 0.0315 0.066872 0.0525 0.0853125 ;
  RECT 0.0315 0.0853125 0.0525 0.139781 ;
  RECT 0.0525 0.066872 0.326813 0.0853125 ;
  RECT 0.326813 0.066872 0.345187 0.0853125 ;
  RECT 0.326813 0.0853125 0.345187 0.139781 ;
  RECT 0.326813 0.139781 0.345187 0.141094 ;
  RECT 0.0958125 0.418687 0.351095 0.437063 ;
  END
END OAI21_X2

MACRO OAI22_X1
  CLASS core ;
  FOREIGN OAI22_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.130594 0.177187 0.378 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.242812 0.183094 0.261188 0.378 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.126 0.135187 0.336 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0315 0.126 0.0525 0.378 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0924655 0.418687 0.200812 0.437063 ;
  RECT 0.200812 0.119437 0.219187 0.418687 ;
  RECT 0.200812 0.418687 0.219187 0.437063 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.261188 0.522375 ;
  RECT 0.261188 0.485625 0.300563 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.300563 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0328125 0.066281 0.242812 0.0859685 ;
  RECT 0.242812 0.066281 0.261188 0.0859685 ;
  RECT 0.242812 0.0859685 0.261188 0.138469 ;
      LAYER M1 ;
  RECT 0.0328125 0.066281 0.242812 0.0859685 ;
  RECT 0.242812 0.066281 0.261188 0.0859685 ;
  RECT 0.242812 0.0859685 0.261188 0.138469 ;
  END
END OAI22_X1

MACRO OAI22_X2
  CLASS core ;
  FOREIGN OAI22_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.504 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.284813 0.168 0.303187 0.183094 ;
  RECT 0.284813 0.183094 0.303187 0.305812 ;
  RECT 0.284813 0.305812 0.303187 0.324188 ;
  RECT 0.303187 0.305812 0.452748 0.324188 ;
  RECT 0.452748 0.183094 0.471187 0.305812 ;
  RECT 0.452748 0.305812 0.471187 0.324188 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.368812 0.168 0.387188 0.261188 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.200812 0.158812 0.219187 0.318937 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.158812 0.093122 0.336 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.253312 0.177187 0.347813 ;
  RECT 0.158812 0.347813 0.177187 0.366187 ;
  RECT 0.177187 0.347813 0.242812 0.366187 ;
  RECT 0.242812 0.110906 0.261188 0.129281 ;
  RECT 0.242812 0.129281 0.261188 0.182437 ;
  RECT 0.242812 0.182437 0.261188 0.253312 ;
  RECT 0.242812 0.253312 0.261188 0.347813 ;
  RECT 0.242812 0.347813 0.261188 0.366187 ;
  RECT 0.261188 0.110906 0.410813 0.129281 ;
  RECT 0.261188 0.347813 0.410813 0.366187 ;
  RECT 0.410813 0.110906 0.429187 0.129281 ;
  RECT 0.410813 0.129281 0.429187 0.182437 ;
  RECT 0.410813 0.347813 0.429187 0.366187 ;
  RECT 0.429187 0.347813 0.452748 0.366187 ;
  RECT 0.452748 0.347813 0.471187 0.366187 ;
  RECT 0.452748 0.366187 0.471187 0.441 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.237562 0.522375 ;
  RECT 0.237562 0.485625 0.429187 0.522375 ;
  RECT 0.429187 0.485625 0.471187 0.522375 ;
  RECT 0.471187 0.485625 0.510565 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.510565 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.263813 0.396375 0.410813 0.417375 ;
  RECT 0.410813 0.396375 0.429187 0.417375 ;
  RECT 0.410813 0.417375 0.429187 0.456685 ;
  RECT 0.0269062 0.064969 0.452748 0.0872815 ;
  RECT 0.452748 0.064969 0.471187 0.0872815 ;
  RECT 0.452748 0.0872815 0.471187 0.138469 ;
  RECT 0.0328125 0.401625 0.237562 0.439688 ;
      LAYER M1 ;
  RECT 0.263813 0.396375 0.410813 0.417375 ;
  RECT 0.410813 0.396375 0.429187 0.417375 ;
  RECT 0.410813 0.417375 0.429187 0.456685 ;
  RECT 0.0269062 0.064969 0.452748 0.0872815 ;
  RECT 0.452748 0.064969 0.471187 0.0872815 ;
  RECT 0.452748 0.0872815 0.471187 0.138469 ;
  RECT 0.0328125 0.401625 0.237562 0.439688 ;
  END
END OAI22_X2

MACRO OR2_X1
  CLASS core ;
  FOREIGN OR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.252 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.063 0.135187 0.336 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.159469 0.0511875 0.420655 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.200812 0.0748125 0.219187 0.42 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.177187 0.522375 ;
  RECT 0.177187 0.485625 0.258562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.258562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0748125 0.0853125 0.093122 0.2205 ;
  RECT 0.0748125 0.2205 0.093122 0.364875 ;
  RECT 0.0748125 0.364875 0.093122 0.38325 ;
  RECT 0.093122 0.364875 0.158812 0.38325 ;
  RECT 0.158812 0.2205 0.177187 0.364875 ;
  RECT 0.158812 0.364875 0.177187 0.38325 ;
      LAYER M1 ;
  RECT 0.0748125 0.0853125 0.093122 0.2205 ;
  RECT 0.0748125 0.2205 0.093122 0.364875 ;
  RECT 0.0748125 0.364875 0.093122 0.38325 ;
  RECT 0.093122 0.364875 0.158812 0.38325 ;
  RECT 0.158812 0.2205 0.177187 0.364875 ;
  RECT 0.158812 0.364875 0.177187 0.38325 ;
  END
END OR2_X1

MACRO OR2_X2
  CLASS core ;
  FOREIGN OR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.294 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.158812 0.093122 0.336 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.168 0.0511875 0.336 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.198187 0.042 0.200812 0.0885935 ;
  RECT 0.198187 0.418687 0.200812 0.462 ;
  RECT 0.200812 0.042 0.219187 0.0885935 ;
  RECT 0.200812 0.0885935 0.219187 0.418687 ;
  RECT 0.200812 0.418687 0.219187 0.462 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.177187 0.522375 ;
  RECT 0.177187 0.485625 0.300563 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.300563 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.050531 0.101062 0.0958125 0.123375 ;
  RECT 0.0958125 0.101062 0.158812 0.123375 ;
  RECT 0.0958125 0.380625 0.158812 0.399 ;
  RECT 0.158812 0.101062 0.177187 0.123375 ;
  RECT 0.158812 0.123375 0.177187 0.380625 ;
  RECT 0.158812 0.380625 0.177187 0.399 ;
      LAYER M1 ;
  RECT 0.050531 0.101062 0.0958125 0.123375 ;
  RECT 0.0958125 0.101062 0.158812 0.123375 ;
  RECT 0.0958125 0.380625 0.158812 0.399 ;
  RECT 0.158812 0.101062 0.177187 0.123375 ;
  RECT 0.158812 0.123375 0.177187 0.380625 ;
  RECT 0.158812 0.380625 0.177187 0.399 ;
  END
END OR2_X2

MACRO OR3_X1
  CLASS core ;
  FOREIGN OR3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.336 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.200812 0.126 0.219187 0.378 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.1155 0.126 0.1365 0.378 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0295312 0.126 0.054469 0.378 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.284813 0.0748125 0.303187 0.429187 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.153562 0.522375 ;
  RECT 0.153562 0.485625 0.261188 0.522375 ;
  RECT 0.261188 0.485625 0.342562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.342562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0354375 0.0715315 0.182437 0.089906 ;
  RECT 0.182437 0.0715315 0.242812 0.089906 ;
  RECT 0.182437 0.414095 0.242812 0.441655 ;
  RECT 0.242812 0.0715315 0.261188 0.089906 ;
  RECT 0.242812 0.089906 0.261188 0.414095 ;
  RECT 0.242812 0.414095 0.261188 0.441655 ;
  RECT 0.056372 0.417375 0.153562 0.438375 ;
      LAYER M1 ;
  RECT 0.0354375 0.0715315 0.182437 0.089906 ;
  RECT 0.182437 0.0715315 0.242812 0.089906 ;
  RECT 0.182437 0.414095 0.242812 0.441655 ;
  RECT 0.242812 0.0715315 0.261188 0.089906 ;
  RECT 0.242812 0.089906 0.261188 0.414095 ;
  RECT 0.242812 0.414095 0.261188 0.441655 ;
  RECT 0.056372 0.417375 0.153562 0.438375 ;
  END
END OR3_X1

MACRO OR3_X2
  CLASS core ;
  FOREIGN OR3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.336 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.167344 0.093122 0.294 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.168 0.0511875 0.345187 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.151594 0.177187 0.294 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.240187 0.042 0.242812 0.0853125 ;
  RECT 0.240187 0.417375 0.242812 0.462 ;
  RECT 0.242812 0.042 0.261188 0.0853125 ;
  RECT 0.242812 0.0853125 0.261188 0.417375 ;
  RECT 0.242812 0.417375 0.261188 0.462 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.198187 0.522375 ;
  RECT 0.198187 0.485625 0.219187 0.522375 ;
  RECT 0.219187 0.485625 0.342562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.342562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0328125 0.375965 0.0511875 0.39572 ;
  RECT 0.0328125 0.39572 0.0511875 0.450188 ;
  RECT 0.0511875 0.375965 0.198187 0.39572 ;
  RECT 0.039375 0.101719 0.0924655 0.122719 ;
  RECT 0.0924655 0.101719 0.200812 0.122719 ;
  RECT 0.0924655 0.331405 0.200812 0.352405 ;
  RECT 0.200812 0.101719 0.219187 0.122719 ;
  RECT 0.200812 0.122719 0.219187 0.331405 ;
  RECT 0.200812 0.331405 0.219187 0.352405 ;
      LAYER M1 ;
  RECT 0.0328125 0.375965 0.0511875 0.39572 ;
  RECT 0.0328125 0.39572 0.0511875 0.450188 ;
  RECT 0.0511875 0.375965 0.198187 0.39572 ;
  RECT 0.039375 0.101719 0.0924655 0.122719 ;
  RECT 0.0924655 0.101719 0.200812 0.122719 ;
  RECT 0.0924655 0.331405 0.200812 0.352405 ;
  RECT 0.200812 0.101719 0.219187 0.122719 ;
  RECT 0.200812 0.122719 0.219187 0.331405 ;
  RECT 0.200812 0.331405 0.219187 0.352405 ;
  END
END OR3_X2

MACRO OR4_X1
  CLASS core ;
  FOREIGN OR4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.378 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.242812 0.126 0.261188 0.378 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.1575 0.126 0.1785 0.378 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.129937 0.093122 0.378 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.126 0.0511875 0.378 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.326813 0.0748125 0.345187 0.42 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.195562 0.522375 ;
  RECT 0.195562 0.485625 0.303187 0.522375 ;
  RECT 0.303187 0.485625 0.384562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.384562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0354375 0.066872 0.221812 0.0853125 ;
  RECT 0.221812 0.066872 0.284813 0.0853125 ;
  RECT 0.221812 0.413438 0.284813 0.434437 ;
  RECT 0.284813 0.066872 0.303187 0.0853125 ;
  RECT 0.284813 0.0853125 0.303187 0.413438 ;
  RECT 0.284813 0.413438 0.303187 0.434437 ;
  RECT 0.0958125 0.404905 0.195562 0.429845 ;
      LAYER M1 ;
  RECT 0.0354375 0.066872 0.221812 0.0853125 ;
  RECT 0.221812 0.066872 0.284813 0.0853125 ;
  RECT 0.221812 0.413438 0.284813 0.434437 ;
  RECT 0.284813 0.066872 0.303187 0.0853125 ;
  RECT 0.284813 0.0853125 0.303187 0.413438 ;
  RECT 0.284813 0.413438 0.303187 0.434437 ;
  RECT 0.0958125 0.404905 0.195562 0.429845 ;
  END
END OR4_X1

MACRO OR4_X2
  CLASS core ;
  FOREIGN OR4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.42 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.200812 0.126 0.219187 0.347813 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.158812 0.139781 0.177187 0.378 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.139781 0.093122 0.378 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.125344 0.0511875 0.378 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.3255 0.084 0.3465 0.462 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.198187 0.522375 ;
  RECT 0.198187 0.485625 0.301875 0.522375 ;
  RECT 0.301875 0.485625 0.426563 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.426563 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0958125 0.408845 0.198187 0.446905 ;
  RECT 0.0354375 0.057028 0.224437 0.095156 ;
  RECT 0.224437 0.057028 0.2835 0.095156 ;
  RECT 0.224437 0.372685 0.2835 0.4095 ;
  RECT 0.2835 0.057028 0.301875 0.095156 ;
  RECT 0.2835 0.095156 0.301875 0.372685 ;
  RECT 0.2835 0.372685 0.301875 0.4095 ;
      LAYER M1 ;
  RECT 0.0958125 0.408845 0.198187 0.446905 ;
  RECT 0.0354375 0.057028 0.224437 0.095156 ;
  RECT 0.224437 0.057028 0.2835 0.095156 ;
  RECT 0.224437 0.372685 0.2835 0.4095 ;
  RECT 0.2835 0.057028 0.301875 0.095156 ;
  RECT 0.2835 0.095156 0.301875 0.372685 ;
  RECT 0.2835 0.372685 0.301875 0.4095 ;
  END
END OR4_X2

MACRO SDFFRNQ_X1
  CLASS core ;
  FOREIGN SDFFRNQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 1.26 BY 0.504 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.326813 0.238219 0.33797 0.3465 ;
  RECT 0.33797 0.238219 0.345187 0.3465 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
  RECT 0.63328 0.221812 0.954185 0.240187 ;
  RECT 0.954185 0.221812 1.04475 0.240187 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.200812 0.244125 0.219187 0.37531 ;
  RECT 0.200812 0.37531 0.219187 0.39375 ;
  RECT 0.219187 0.37531 0.33797 0.39375 ;
  RECT 0.33797 0.37531 0.368812 0.39375 ;
  RECT 0.368812 0.206062 0.387188 0.244125 ;
  RECT 0.368812 0.244125 0.387188 0.37531 ;
  RECT 0.368812 0.37531 0.387188 0.39375 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.242812 0.238219 0.261188 0.336 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.181125 0.0511875 0.350438 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 1.2075 0.042 1.2285 0.462 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.093122 0.522375 ;
  RECT 0.093122 0.485625 0.135187 0.522375 ;
  RECT 0.135187 0.485625 0.494812 0.522375 ;
  RECT 0.494812 0.485625 0.51319 0.522375 ;
  RECT 0.51319 0.485625 0.69956 0.522375 ;
  RECT 0.69956 0.485625 0.933185 0.522375 ;
  RECT 0.933185 0.485625 0.97781 0.522375 ;
  RECT 0.97781 0.485625 1.14319 0.522375 ;
  RECT 1.14319 0.485625 1.26656 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 1.26656 0.018375 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
  RECT 0.0958125 0.347813 0.87019 0.366187 ;
  RECT 0.473813 0.263813 0.735655 0.282187 ;
  RECT 0.0538125 0.179812 0.954185 0.198187 ;
      LAYER MINT1 ;
  RECT 0.0958125 0.347813 0.87019 0.366187 ;
  RECT 0.473813 0.263813 0.735655 0.282187 ;
  RECT 0.0538125 0.179812 0.954185 0.198187 ;
      LAYER M1 ;
  RECT 0.0295312 0.063 0.054469 0.133809 ;
  RECT 0.0295312 0.133809 0.054469 0.15225 ;
  RECT 0.0295312 0.396375 0.054469 0.41475 ;
  RECT 0.0295312 0.41475 0.054469 0.451435 ;
  RECT 0.054469 0.133809 0.0748125 0.15225 ;
  RECT 0.054469 0.396375 0.0748125 0.41475 ;
  RECT 0.0748125 0.133809 0.093122 0.15225 ;
  RECT 0.0748125 0.15225 0.093122 0.396375 ;
  RECT 0.0748125 0.396375 0.093122 0.41475 ;
  RECT 0.158812 0.063 0.177187 0.175219 ;
  RECT 0.158812 0.175219 0.177187 0.193594 ;
  RECT 0.158812 0.193594 0.177187 0.441 ;
  RECT 0.177187 0.175219 0.33797 0.193594 ;
  RECT 0.221812 0.12075 0.410813 0.139125 ;
  RECT 0.410813 0.12075 0.429187 0.139125 ;
  RECT 0.410813 0.139125 0.429187 0.181125 ;
  RECT 0.25725 0.417375 0.494812 0.438375 ;
  RECT 0.494812 0.162094 0.51319 0.358312 ;
  RECT 0.305812 0.066872 0.576185 0.0853125 ;
  RECT 0.69628 0.1575 0.72056 0.292687 ;
  RECT 0.788815 0.112219 0.807185 0.335345 ;
  RECT 0.95681 0.0958125 0.97781 0.457998 ;
  RECT 0.76453 0.405562 0.87281 0.423938 ;
  RECT 0.87281 0.042 0.89119 0.060375 ;
  RECT 0.87281 0.060375 0.89119 0.240187 ;
  RECT 0.87281 0.240187 0.89119 0.405562 ;
  RECT 0.87281 0.405562 0.89119 0.423938 ;
  RECT 0.89119 0.042 1.05459 0.060375 ;
  RECT 1.05459 0.042 1.07297 0.060375 ;
  RECT 1.05459 0.060375 1.07297 0.240187 ;
  RECT 1.01981 0.301875 1.03819 0.4095 ;
  RECT 1.01981 0.4095 1.03819 0.44625 ;
  RECT 1.03819 0.4095 1.12481 0.44625 ;
  RECT 1.12481 0.04725 1.14319 0.301875 ;
  RECT 1.12481 0.301875 1.14319 0.4095 ;
  RECT 1.12481 0.4095 1.14319 0.44625 ;
  RECT 0.116812 0.082031 0.135187 0.376688 ;
  RECT 0.452748 0.25397 0.471187 0.387188 ;
  RECT 0.53675 0.168656 0.557815 0.30778 ;
  RECT 0.452748 0.108937 0.471187 0.127312 ;
  RECT 0.452748 0.127312 0.471187 0.181125 ;
  RECT 0.471187 0.108937 0.61819 0.127312 ;
  RECT 0.650345 0.158812 0.672655 0.276938 ;
  RECT 0.518435 0.417375 0.69956 0.438375 ;
  RECT 0.59325 0.179812 0.611625 0.321562 ;
  RECT 0.59325 0.321562 0.611625 0.339938 ;
  RECT 0.611625 0.321562 0.744125 0.339938 ;
  RECT 0.744125 0.0538125 0.76519 0.179812 ;
  RECT 0.744125 0.179812 0.76519 0.321562 ;
  RECT 0.744125 0.321562 0.76519 0.339938 ;
  RECT 0.83081 0.116812 0.849185 0.376688 ;
  RECT 0.91475 0.116812 0.933185 0.324188 ;
  RECT 1.00537 0.101062 1.03097 0.273 ;
      LAYER V1 ;
  RECT 0.0748125 0.179812 0.093122 0.198187 ;
  RECT 0.116812 0.347813 0.135187 0.366187 ;
  RECT 0.452748 0.347813 0.471187 0.366187 ;
  RECT 0.494812 0.263813 0.51319 0.282187 ;
  RECT 0.53675 0.179812 0.555185 0.198187 ;
  RECT 0.65428 0.221812 0.672655 0.240187 ;
  RECT 0.69628 0.263813 0.714655 0.282187 ;
  RECT 0.788815 0.179812 0.807185 0.198187 ;
  RECT 0.83081 0.347813 0.849185 0.366187 ;
  RECT 0.91475 0.179812 0.933185 0.198187 ;
  RECT 1.00537 0.221812 1.02375 0.240187 ;
      LAYER M1 ;
  RECT 0.0295312 0.063 0.054469 0.133809 ;
  RECT 0.0295312 0.133809 0.054469 0.15225 ;
  RECT 0.0295312 0.396375 0.054469 0.41475 ;
  RECT 0.0295312 0.41475 0.054469 0.451435 ;
  RECT 0.054469 0.133809 0.0748125 0.15225 ;
  RECT 0.054469 0.396375 0.0748125 0.41475 ;
  RECT 0.0748125 0.133809 0.093122 0.15225 ;
  RECT 0.0748125 0.15225 0.093122 0.396375 ;
  RECT 0.0748125 0.396375 0.093122 0.41475 ;
  RECT 0.158812 0.063 0.177187 0.175219 ;
  RECT 0.158812 0.175219 0.177187 0.193594 ;
  RECT 0.158812 0.193594 0.177187 0.441 ;
  RECT 0.177187 0.175219 0.33797 0.193594 ;
  RECT 0.221812 0.12075 0.410813 0.139125 ;
  RECT 0.410813 0.12075 0.429187 0.139125 ;
  RECT 0.410813 0.139125 0.429187 0.181125 ;
  RECT 0.25725 0.417375 0.494812 0.438375 ;
  RECT 0.494812 0.162094 0.51319 0.358312 ;
  RECT 0.305812 0.066872 0.576185 0.0853125 ;
  RECT 0.69628 0.1575 0.72056 0.292687 ;
  RECT 0.788815 0.112219 0.807185 0.335345 ;
  RECT 0.95681 0.0958125 0.97781 0.457998 ;
  RECT 0.76453 0.405562 0.87281 0.423938 ;
  RECT 0.87281 0.042 0.89119 0.060375 ;
  RECT 0.87281 0.060375 0.89119 0.240187 ;
  RECT 0.87281 0.240187 0.89119 0.405562 ;
  RECT 0.87281 0.405562 0.89119 0.423938 ;
  RECT 0.89119 0.042 1.05459 0.060375 ;
  RECT 1.05459 0.042 1.07297 0.060375 ;
  RECT 1.05459 0.060375 1.07297 0.240187 ;
  RECT 1.01981 0.301875 1.03819 0.4095 ;
  RECT 1.01981 0.4095 1.03819 0.44625 ;
  RECT 1.03819 0.4095 1.12481 0.44625 ;
  RECT 1.12481 0.04725 1.14319 0.301875 ;
  RECT 1.12481 0.301875 1.14319 0.4095 ;
  RECT 1.12481 0.4095 1.14319 0.44625 ;
  RECT 0.116812 0.082031 0.135187 0.376688 ;
  RECT 0.452748 0.25397 0.471187 0.387188 ;
  RECT 0.53675 0.168656 0.557815 0.30778 ;
  RECT 0.452748 0.108937 0.471187 0.127312 ;
  RECT 0.452748 0.127312 0.471187 0.181125 ;
  RECT 0.471187 0.108937 0.61819 0.127312 ;
  RECT 0.650345 0.158812 0.672655 0.276938 ;
  RECT 0.518435 0.417375 0.69956 0.438375 ;
  RECT 0.59325 0.179812 0.611625 0.321562 ;
  RECT 0.59325 0.321562 0.611625 0.339938 ;
  RECT 0.611625 0.321562 0.744125 0.339938 ;
  RECT 0.744125 0.0538125 0.76519 0.179812 ;
  RECT 0.744125 0.179812 0.76519 0.321562 ;
  RECT 0.744125 0.321562 0.76519 0.339938 ;
  RECT 0.83081 0.116812 0.849185 0.376688 ;
  RECT 0.91475 0.116812 0.933185 0.324188 ;
  RECT 1.00537 0.101062 1.03097 0.273 ;
  END
END SDFFRNQ_X1

MACRO SDFFSNQ_X1
  CLASS core ;
  FOREIGN SDFFSNQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 1.26 BY 0.504 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.326813 0.252 0.334688 0.3465 ;
  RECT 0.334688 0.252 0.345187 0.3465 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.200812 0.244125 0.219187 0.37531 ;
  RECT 0.200812 0.37531 0.219187 0.39375 ;
  RECT 0.219187 0.37531 0.334688 0.39375 ;
  RECT 0.334688 0.37531 0.368812 0.39375 ;
  RECT 0.368812 0.206062 0.387188 0.244125 ;
  RECT 0.368812 0.244125 0.387188 0.37531 ;
  RECT 0.368812 0.37531 0.387188 0.39375 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.242812 0.238219 0.261188 0.336 ;
    END
  END SI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
  RECT 0.628685 0.221812 0.954185 0.240187 ;
  RECT 0.954185 0.221812 1.04081 0.240187 ;
    END
  END SN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.1785 0.0511875 0.336 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 1.2075 0.042 1.2285 0.462 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.093122 0.522375 ;
  RECT 0.093122 0.485625 0.135187 0.522375 ;
  RECT 0.135187 0.485625 0.489563 0.522375 ;
  RECT 0.489563 0.485625 0.51319 0.522375 ;
  RECT 0.51319 0.485625 0.56569 0.522375 ;
  RECT 0.56569 0.485625 1.08019 0.522375 ;
  RECT 1.08019 0.485625 1.14319 0.522375 ;
  RECT 1.14319 0.485625 1.26656 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 1.26656 0.018375 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
  RECT 0.0958125 0.347813 0.87019 0.366187 ;
  RECT 0.473813 0.263813 0.73106 0.282187 ;
  RECT 0.0538125 0.179812 0.954185 0.198187 ;
      LAYER MINT1 ;
  RECT 0.0958125 0.347813 0.87019 0.366187 ;
  RECT 0.473813 0.263813 0.73106 0.282187 ;
  RECT 0.0538125 0.179812 0.954185 0.198187 ;
      LAYER M1 ;
  RECT 0.0315 0.042 0.0525 0.13125 ;
  RECT 0.0315 0.13125 0.0525 0.149625 ;
  RECT 0.0315 0.396375 0.0525 0.41475 ;
  RECT 0.0315 0.41475 0.0525 0.451435 ;
  RECT 0.0525 0.13125 0.0748125 0.149625 ;
  RECT 0.0525 0.396375 0.0748125 0.41475 ;
  RECT 0.0748125 0.13125 0.093122 0.149625 ;
  RECT 0.0748125 0.149625 0.093122 0.396375 ;
  RECT 0.0748125 0.396375 0.093122 0.41475 ;
  RECT 0.158812 0.0538125 0.177187 0.174562 ;
  RECT 0.158812 0.174562 0.177187 0.193594 ;
  RECT 0.158812 0.193594 0.177187 0.19425 ;
  RECT 0.158812 0.19425 0.177187 0.450188 ;
  RECT 0.177187 0.174562 0.284813 0.193594 ;
  RECT 0.284813 0.174562 0.334688 0.193594 ;
  RECT 0.284813 0.193594 0.334688 0.19425 ;
  RECT 0.221812 0.12075 0.410813 0.139125 ;
  RECT 0.410813 0.12075 0.429187 0.139125 ;
  RECT 0.410813 0.139125 0.429187 0.181125 ;
  RECT 0.25725 0.417375 0.489563 0.438375 ;
  RECT 0.494812 0.156187 0.51319 0.35897 ;
  RECT 0.305812 0.066872 0.576185 0.0853125 ;
  RECT 0.643125 0.211312 0.668065 0.27497 ;
  RECT 0.589315 0.179812 0.60769 0.319595 ;
  RECT 0.589315 0.319595 0.60769 0.33797 ;
  RECT 0.60769 0.319595 0.6615 0.33797 ;
  RECT 0.6615 0.319595 0.6825 0.33797 ;
  RECT 0.6615 0.33797 0.6825 0.462 ;
  RECT 0.6825 0.319595 0.74675 0.33797 ;
  RECT 0.74675 0.0643125 0.76519 0.179812 ;
  RECT 0.74675 0.179812 0.76519 0.319595 ;
  RECT 0.74675 0.319595 0.76519 0.33797 ;
  RECT 0.83081 0.116812 0.849185 0.376688 ;
  RECT 0.91475 0.116812 0.933185 0.263813 ;
  RECT 1.00144 0.12075 1.01981 0.26447 ;
  RECT 0.920065 0.418687 1.08019 0.437063 ;
  RECT 0.116812 0.063 0.135187 0.40622 ;
  RECT 0.429187 0.25397 0.447562 0.376688 ;
  RECT 0.544685 0.168656 0.56569 0.30778 ;
  RECT 0.452748 0.108937 0.471187 0.127312 ;
  RECT 0.452748 0.127312 0.471187 0.181125 ;
  RECT 0.471187 0.108937 0.61819 0.127312 ;
  RECT 0.69169 0.1575 0.716625 0.292687 ;
  RECT 0.788815 0.112219 0.807185 0.251345 ;
  RECT 0.76453 0.405562 0.87281 0.423938 ;
  RECT 0.87281 0.0538125 0.89119 0.0721875 ;
  RECT 0.87281 0.0721875 0.89119 0.240187 ;
  RECT 0.87281 0.240187 0.89119 0.405562 ;
  RECT 0.87281 0.405562 0.89119 0.423938 ;
  RECT 0.89119 0.0538125 1.05459 0.0721875 ;
  RECT 1.05459 0.0538125 1.07953 0.0721875 ;
  RECT 1.05459 0.0721875 1.07953 0.240187 ;
  RECT 0.95944 0.263813 0.97781 0.376688 ;
  RECT 0.95944 0.376688 0.97781 0.395062 ;
  RECT 0.97781 0.376688 1.12481 0.395062 ;
  RECT 1.12481 0.063 1.14319 0.263813 ;
  RECT 1.12481 0.263813 1.14319 0.376688 ;
  RECT 1.12481 0.376688 1.14319 0.395062 ;
      LAYER V1 ;
  RECT 0.0748125 0.179812 0.093122 0.198187 ;
  RECT 0.116812 0.347813 0.135187 0.366187 ;
  RECT 0.429187 0.347813 0.447562 0.366187 ;
  RECT 0.494812 0.263813 0.51319 0.282187 ;
  RECT 0.54731 0.179812 0.56569 0.198187 ;
  RECT 0.649685 0.221812 0.668065 0.240187 ;
  RECT 0.69169 0.263813 0.710065 0.282187 ;
  RECT 0.788815 0.179812 0.807185 0.198187 ;
  RECT 0.83081 0.347813 0.849185 0.366187 ;
  RECT 0.91475 0.179812 0.933185 0.198187 ;
  RECT 1.00144 0.221812 1.01981 0.240187 ;
      LAYER M1 ;
  RECT 0.0315 0.042 0.0525 0.13125 ;
  RECT 0.0315 0.13125 0.0525 0.149625 ;
  RECT 0.0315 0.396375 0.0525 0.41475 ;
  RECT 0.0315 0.41475 0.0525 0.451435 ;
  RECT 0.0525 0.13125 0.0748125 0.149625 ;
  RECT 0.0525 0.396375 0.0748125 0.41475 ;
  RECT 0.0748125 0.13125 0.093122 0.149625 ;
  RECT 0.0748125 0.149625 0.093122 0.396375 ;
  RECT 0.0748125 0.396375 0.093122 0.41475 ;
  RECT 0.158812 0.0538125 0.177187 0.174562 ;
  RECT 0.158812 0.174562 0.177187 0.193594 ;
  RECT 0.158812 0.193594 0.177187 0.19425 ;
  RECT 0.158812 0.19425 0.177187 0.450188 ;
  RECT 0.177187 0.174562 0.284813 0.193594 ;
  RECT 0.284813 0.174562 0.334688 0.193594 ;
  RECT 0.284813 0.193594 0.334688 0.19425 ;
  RECT 0.221812 0.12075 0.410813 0.139125 ;
  RECT 0.410813 0.12075 0.429187 0.139125 ;
  RECT 0.410813 0.139125 0.429187 0.181125 ;
  RECT 0.25725 0.417375 0.489563 0.438375 ;
  RECT 0.494812 0.156187 0.51319 0.35897 ;
  RECT 0.305812 0.066872 0.576185 0.0853125 ;
  RECT 0.643125 0.211312 0.668065 0.27497 ;
  RECT 0.589315 0.179812 0.60769 0.319595 ;
  RECT 0.589315 0.319595 0.60769 0.33797 ;
  RECT 0.60769 0.319595 0.6615 0.33797 ;
  RECT 0.6615 0.319595 0.6825 0.33797 ;
  RECT 0.6615 0.33797 0.6825 0.462 ;
  RECT 0.6825 0.319595 0.74675 0.33797 ;
  RECT 0.74675 0.0643125 0.76519 0.179812 ;
  RECT 0.74675 0.179812 0.76519 0.319595 ;
  RECT 0.74675 0.319595 0.76519 0.33797 ;
  RECT 0.83081 0.116812 0.849185 0.376688 ;
  RECT 0.91475 0.116812 0.933185 0.263813 ;
  RECT 1.00144 0.12075 1.01981 0.26447 ;
  RECT 0.920065 0.418687 1.08019 0.437063 ;
  RECT 0.116812 0.063 0.135187 0.40622 ;
  RECT 0.429187 0.25397 0.447562 0.376688 ;
  RECT 0.544685 0.168656 0.56569 0.30778 ;
  RECT 0.452748 0.108937 0.471187 0.127312 ;
  RECT 0.452748 0.127312 0.471187 0.181125 ;
  RECT 0.471187 0.108937 0.61819 0.127312 ;
  RECT 0.69169 0.1575 0.716625 0.292687 ;
  RECT 0.788815 0.112219 0.807185 0.251345 ;
  RECT 0.76453 0.405562 0.87281 0.423938 ;
  RECT 0.87281 0.0538125 0.89119 0.0721875 ;
  RECT 0.87281 0.0721875 0.89119 0.240187 ;
  RECT 0.87281 0.240187 0.89119 0.405562 ;
  RECT 0.87281 0.405562 0.89119 0.423938 ;
  RECT 0.89119 0.0538125 1.05459 0.0721875 ;
  RECT 1.05459 0.0538125 1.07953 0.0721875 ;
  RECT 1.05459 0.0721875 1.07953 0.240187 ;
  RECT 0.95944 0.263813 0.97781 0.376688 ;
  RECT 0.95944 0.376688 0.97781 0.395062 ;
  RECT 0.97781 0.376688 1.12481 0.395062 ;
  RECT 1.12481 0.063 1.14319 0.263813 ;
  RECT 1.12481 0.263813 1.14319 0.376688 ;
  RECT 1.12481 0.376688 1.14319 0.395062 ;
  END
END SDFFSNQ_X1

MACRO TBUF_X1
  CLASS core ;
  FOREIGN TBUF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.462 BY 0.504 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.252 0.093122 0.322875 ;
  RECT 0.0748125 0.322875 0.093122 0.34125 ;
  RECT 0.093122 0.322875 0.135187 0.34125 ;
  RECT 0.135187 0.322875 0.158812 0.34125 ;
  RECT 0.158812 0.200812 0.177187 0.252 ;
  RECT 0.158812 0.252 0.177187 0.322875 ;
  RECT 0.158812 0.322875 0.177187 0.34125 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.284813 0.242812 0.303187 0.378 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.4095 0.042 0.4305 0.462 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.385875 0.522375 ;
  RECT 0.385875 0.485625 0.468562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.468562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0328125 0.04725 0.0511875 0.20475 ;
  RECT 0.0328125 0.20475 0.0511875 0.223125 ;
  RECT 0.0328125 0.223125 0.0511875 0.274313 ;
  RECT 0.0328125 0.274313 0.0511875 0.450188 ;
  RECT 0.0511875 0.20475 0.116812 0.223125 ;
  RECT 0.116812 0.20475 0.135187 0.223125 ;
  RECT 0.116812 0.223125 0.135187 0.274313 ;
  RECT 0.0958125 0.376688 0.132562 0.395062 ;
  RECT 0.132562 0.066872 0.150937 0.0853125 ;
  RECT 0.132562 0.0853125 0.150937 0.150937 ;
  RECT 0.132562 0.150937 0.150937 0.169312 ;
  RECT 0.132562 0.376688 0.150937 0.395062 ;
  RECT 0.150937 0.066872 0.200812 0.0853125 ;
  RECT 0.150937 0.150937 0.200812 0.169312 ;
  RECT 0.150937 0.376688 0.200812 0.395062 ;
  RECT 0.200812 0.066872 0.219187 0.0853125 ;
  RECT 0.200812 0.150937 0.219187 0.169312 ;
  RECT 0.200812 0.169312 0.219187 0.206062 ;
  RECT 0.200812 0.206062 0.219187 0.376688 ;
  RECT 0.200812 0.376688 0.219187 0.395062 ;
  RECT 0.219187 0.066872 0.334688 0.0853125 ;
  RECT 0.334688 0.066872 0.355687 0.0853125 ;
  RECT 0.334688 0.0853125 0.355687 0.150937 ;
  RECT 0.334688 0.150937 0.355687 0.169312 ;
  RECT 0.334688 0.169312 0.355687 0.206062 ;
  RECT 0.0958125 0.418687 0.179812 0.437063 ;
  RECT 0.179812 0.108937 0.242812 0.127312 ;
  RECT 0.179812 0.418687 0.242812 0.437063 ;
  RECT 0.242812 0.108937 0.261188 0.127312 ;
  RECT 0.242812 0.127312 0.261188 0.24675 ;
  RECT 0.242812 0.24675 0.261188 0.418687 ;
  RECT 0.242812 0.418687 0.261188 0.437063 ;
  RECT 0.261188 0.418687 0.3675 0.437063 ;
  RECT 0.3675 0.24675 0.385875 0.418687 ;
  RECT 0.3675 0.418687 0.385875 0.437063 ;
      LAYER M1 ;
  RECT 0.0328125 0.04725 0.0511875 0.20475 ;
  RECT 0.0328125 0.20475 0.0511875 0.223125 ;
  RECT 0.0328125 0.223125 0.0511875 0.274313 ;
  RECT 0.0328125 0.274313 0.0511875 0.450188 ;
  RECT 0.0511875 0.20475 0.116812 0.223125 ;
  RECT 0.116812 0.20475 0.135187 0.223125 ;
  RECT 0.116812 0.223125 0.135187 0.274313 ;
  RECT 0.0958125 0.376688 0.132562 0.395062 ;
  RECT 0.132562 0.066872 0.150937 0.0853125 ;
  RECT 0.132562 0.0853125 0.150937 0.150937 ;
  RECT 0.132562 0.150937 0.150937 0.169312 ;
  RECT 0.132562 0.376688 0.150937 0.395062 ;
  RECT 0.150937 0.066872 0.200812 0.0853125 ;
  RECT 0.150937 0.150937 0.200812 0.169312 ;
  RECT 0.150937 0.376688 0.200812 0.395062 ;
  RECT 0.200812 0.066872 0.219187 0.0853125 ;
  RECT 0.200812 0.150937 0.219187 0.169312 ;
  RECT 0.200812 0.169312 0.219187 0.206062 ;
  RECT 0.200812 0.206062 0.219187 0.376688 ;
  RECT 0.200812 0.376688 0.219187 0.395062 ;
  RECT 0.219187 0.066872 0.334688 0.0853125 ;
  RECT 0.334688 0.066872 0.355687 0.0853125 ;
  RECT 0.334688 0.0853125 0.355687 0.150937 ;
  RECT 0.334688 0.150937 0.355687 0.169312 ;
  RECT 0.334688 0.169312 0.355687 0.206062 ;
  RECT 0.0958125 0.418687 0.179812 0.437063 ;
  RECT 0.179812 0.108937 0.242812 0.127312 ;
  RECT 0.179812 0.418687 0.242812 0.437063 ;
  RECT 0.242812 0.108937 0.261188 0.127312 ;
  RECT 0.242812 0.127312 0.261188 0.24675 ;
  RECT 0.242812 0.24675 0.261188 0.418687 ;
  RECT 0.242812 0.418687 0.261188 0.437063 ;
  RECT 0.261188 0.418687 0.3675 0.437063 ;
  RECT 0.3675 0.24675 0.385875 0.418687 ;
  RECT 0.3675 0.418687 0.385875 0.437063 ;
  END
END TBUF_X1

MACRO TBUF_X2
  CLASS core ;
  FOREIGN TBUF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.504 BY 0.504 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.252 0.093122 0.33075 ;
  RECT 0.0748125 0.33075 0.093122 0.349125 ;
  RECT 0.093122 0.33075 0.135187 0.349125 ;
  RECT 0.135187 0.33075 0.158812 0.349125 ;
  RECT 0.158812 0.200812 0.177187 0.252 ;
  RECT 0.158812 0.252 0.177187 0.33075 ;
  RECT 0.158812 0.33075 0.177187 0.349125 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.284813 0.250688 0.303187 0.378 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.4095 0.0459375 0.4305 0.456685 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.347813 0.522375 ;
  RECT 0.347813 0.485625 0.510565 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.510565 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0328125 0.04725 0.0511875 0.20475 ;
  RECT 0.0328125 0.20475 0.0511875 0.223125 ;
  RECT 0.0328125 0.223125 0.0511875 0.265125 ;
  RECT 0.0328125 0.265125 0.0511875 0.401625 ;
  RECT 0.0511875 0.20475 0.116812 0.223125 ;
  RECT 0.116812 0.20475 0.135187 0.223125 ;
  RECT 0.116812 0.223125 0.135187 0.265125 ;
  RECT 0.0958125 0.372685 0.132562 0.395062 ;
  RECT 0.132562 0.066872 0.150937 0.0853125 ;
  RECT 0.132562 0.0853125 0.150937 0.150937 ;
  RECT 0.132562 0.150937 0.150937 0.169312 ;
  RECT 0.132562 0.372685 0.150937 0.395062 ;
  RECT 0.150937 0.066872 0.200812 0.0853125 ;
  RECT 0.150937 0.150937 0.200812 0.169312 ;
  RECT 0.150937 0.372685 0.200812 0.395062 ;
  RECT 0.200812 0.066872 0.219187 0.0853125 ;
  RECT 0.200812 0.150937 0.219187 0.169312 ;
  RECT 0.200812 0.169312 0.219187 0.206062 ;
  RECT 0.200812 0.206062 0.219187 0.372685 ;
  RECT 0.200812 0.372685 0.219187 0.395062 ;
  RECT 0.219187 0.066872 0.316312 0.0853125 ;
  RECT 0.316312 0.066872 0.337313 0.0853125 ;
  RECT 0.316312 0.0853125 0.337313 0.150937 ;
  RECT 0.316312 0.150937 0.337313 0.169312 ;
  RECT 0.316312 0.169312 0.337313 0.206062 ;
  RECT 0.0958125 0.418687 0.179812 0.437063 ;
  RECT 0.179812 0.108937 0.242812 0.127312 ;
  RECT 0.179812 0.418687 0.242812 0.437063 ;
  RECT 0.242812 0.108937 0.261188 0.127312 ;
  RECT 0.242812 0.127312 0.261188 0.29072 ;
  RECT 0.242812 0.29072 0.261188 0.418687 ;
  RECT 0.242812 0.418687 0.261188 0.437063 ;
  RECT 0.261188 0.418687 0.326813 0.437063 ;
  RECT 0.326813 0.29072 0.347813 0.418687 ;
  RECT 0.326813 0.418687 0.347813 0.437063 ;
      LAYER M1 ;
  RECT 0.0328125 0.04725 0.0511875 0.20475 ;
  RECT 0.0328125 0.20475 0.0511875 0.223125 ;
  RECT 0.0328125 0.223125 0.0511875 0.265125 ;
  RECT 0.0328125 0.265125 0.0511875 0.401625 ;
  RECT 0.0511875 0.20475 0.116812 0.223125 ;
  RECT 0.116812 0.20475 0.135187 0.223125 ;
  RECT 0.116812 0.223125 0.135187 0.265125 ;
  RECT 0.0958125 0.372685 0.132562 0.395062 ;
  RECT 0.132562 0.066872 0.150937 0.0853125 ;
  RECT 0.132562 0.0853125 0.150937 0.150937 ;
  RECT 0.132562 0.150937 0.150937 0.169312 ;
  RECT 0.132562 0.372685 0.150937 0.395062 ;
  RECT 0.150937 0.066872 0.200812 0.0853125 ;
  RECT 0.150937 0.150937 0.200812 0.169312 ;
  RECT 0.150937 0.372685 0.200812 0.395062 ;
  RECT 0.200812 0.066872 0.219187 0.0853125 ;
  RECT 0.200812 0.150937 0.219187 0.169312 ;
  RECT 0.200812 0.169312 0.219187 0.206062 ;
  RECT 0.200812 0.206062 0.219187 0.372685 ;
  RECT 0.200812 0.372685 0.219187 0.395062 ;
  RECT 0.219187 0.066872 0.316312 0.0853125 ;
  RECT 0.316312 0.066872 0.337313 0.0853125 ;
  RECT 0.316312 0.0853125 0.337313 0.150937 ;
  RECT 0.316312 0.150937 0.337313 0.169312 ;
  RECT 0.316312 0.169312 0.337313 0.206062 ;
  RECT 0.0958125 0.418687 0.179812 0.437063 ;
  RECT 0.179812 0.108937 0.242812 0.127312 ;
  RECT 0.179812 0.418687 0.242812 0.437063 ;
  RECT 0.242812 0.108937 0.261188 0.127312 ;
  RECT 0.242812 0.127312 0.261188 0.29072 ;
  RECT 0.242812 0.29072 0.261188 0.418687 ;
  RECT 0.242812 0.418687 0.261188 0.437063 ;
  RECT 0.261188 0.418687 0.326813 0.437063 ;
  RECT 0.326813 0.29072 0.347813 0.418687 ;
  RECT 0.326813 0.418687 0.347813 0.437063 ;
  END
END TBUF_X2

MACRO TBUF_X4
  CLASS core ;
  FOREIGN TBUF_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.63 BY 0.504 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.252 0.093122 0.317625 ;
  RECT 0.0748125 0.317625 0.093122 0.336 ;
  RECT 0.093122 0.317625 0.135187 0.336 ;
  RECT 0.135187 0.317625 0.158812 0.336 ;
  RECT 0.158812 0.200812 0.177187 0.252 ;
  RECT 0.158812 0.252 0.177187 0.317625 ;
  RECT 0.158812 0.317625 0.177187 0.336 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.284813 0.226997 0.303187 0.389813 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.451435 0.042 0.4725 0.147 ;
  RECT 0.451435 0.147 0.4725 0.168 ;
  RECT 0.451435 0.336 0.4725 0.354375 ;
  RECT 0.451435 0.354375 0.4725 0.374652 ;
  RECT 0.451435 0.374652 0.4725 0.462 ;
  RECT 0.4725 0.147 0.533465 0.168 ;
  RECT 0.4725 0.336 0.533465 0.354375 ;
  RECT 0.533465 0.042 0.53412 0.147 ;
  RECT 0.533465 0.147 0.53412 0.168 ;
  RECT 0.533465 0.336 0.53412 0.354375 ;
  RECT 0.53412 0.042 0.535435 0.147 ;
  RECT 0.53412 0.147 0.535435 0.168 ;
  RECT 0.53412 0.336 0.535435 0.354375 ;
  RECT 0.535435 0.042 0.549935 0.147 ;
  RECT 0.535435 0.147 0.549935 0.168 ;
  RECT 0.535435 0.336 0.549935 0.354375 ;
  RECT 0.535435 0.354375 0.549935 0.374652 ;
  RECT 0.535435 0.374652 0.549935 0.462 ;
  RECT 0.549935 0.042 0.5565 0.147 ;
  RECT 0.549935 0.147 0.5565 0.168 ;
  RECT 0.549935 0.336 0.5565 0.354375 ;
  RECT 0.549935 0.354375 0.5565 0.374652 ;
  RECT 0.549935 0.374652 0.5565 0.462 ;
  RECT 0.5565 0.042 0.55847 0.147 ;
  RECT 0.5565 0.147 0.55847 0.168 ;
  RECT 0.5565 0.336 0.55847 0.354375 ;
  RECT 0.5565 0.354375 0.55847 0.374652 ;
  RECT 0.55847 0.147 0.57881 0.168 ;
  RECT 0.55847 0.336 0.57881 0.354375 ;
  RECT 0.55847 0.354375 0.57881 0.374652 ;
  RECT 0.57881 0.147 0.597185 0.168 ;
  RECT 0.57881 0.168 0.597185 0.336 ;
  RECT 0.57881 0.336 0.597185 0.354375 ;
  RECT 0.57881 0.354375 0.597185 0.374652 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.53412 0.522375 ;
  RECT 0.53412 0.485625 0.549935 0.522375 ;
  RECT 0.549935 0.485625 0.636565 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.636565 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0538125 0.418687 0.179812 0.437063 ;
  RECT 0.179812 0.108937 0.242812 0.127312 ;
  RECT 0.179812 0.418687 0.242812 0.437063 ;
  RECT 0.242812 0.108937 0.261188 0.127312 ;
  RECT 0.242812 0.127312 0.261188 0.254625 ;
  RECT 0.242812 0.254625 0.261188 0.271688 ;
  RECT 0.242812 0.271688 0.261188 0.300563 ;
  RECT 0.242812 0.300563 0.261188 0.418687 ;
  RECT 0.242812 0.418687 0.261188 0.437063 ;
  RECT 0.261188 0.418687 0.345187 0.437063 ;
  RECT 0.345187 0.254625 0.381937 0.271688 ;
  RECT 0.345187 0.271688 0.381937 0.300563 ;
  RECT 0.345187 0.300563 0.381937 0.418687 ;
  RECT 0.345187 0.418687 0.381937 0.437063 ;
  RECT 0.381937 0.271688 0.53412 0.300563 ;
  RECT 0.0328125 0.063 0.0511875 0.20475 ;
  RECT 0.0328125 0.20475 0.0511875 0.223125 ;
  RECT 0.0328125 0.223125 0.0511875 0.265125 ;
  RECT 0.0328125 0.265125 0.0511875 0.389813 ;
  RECT 0.0511875 0.20475 0.116812 0.223125 ;
  RECT 0.116812 0.20475 0.135187 0.223125 ;
  RECT 0.116812 0.223125 0.135187 0.265125 ;
  RECT 0.0958125 0.372685 0.132562 0.395062 ;
  RECT 0.132562 0.066872 0.150937 0.0853125 ;
  RECT 0.132562 0.0853125 0.150937 0.150937 ;
  RECT 0.132562 0.150937 0.150937 0.169312 ;
  RECT 0.132562 0.372685 0.150937 0.395062 ;
  RECT 0.150937 0.066872 0.200812 0.0853125 ;
  RECT 0.150937 0.150937 0.200812 0.169312 ;
  RECT 0.150937 0.372685 0.200812 0.395062 ;
  RECT 0.200812 0.066872 0.219187 0.0853125 ;
  RECT 0.200812 0.150937 0.219187 0.169312 ;
  RECT 0.200812 0.169312 0.219187 0.191625 ;
  RECT 0.200812 0.191625 0.219187 0.21 ;
  RECT 0.200812 0.21 0.219187 0.231 ;
  RECT 0.200812 0.231 0.219187 0.372685 ;
  RECT 0.200812 0.372685 0.219187 0.395062 ;
  RECT 0.219187 0.066872 0.345187 0.0853125 ;
  RECT 0.345187 0.066872 0.381937 0.0853125 ;
  RECT 0.345187 0.0853125 0.381937 0.150937 ;
  RECT 0.345187 0.150937 0.381937 0.169312 ;
  RECT 0.345187 0.169312 0.381937 0.191625 ;
  RECT 0.345187 0.191625 0.381937 0.21 ;
  RECT 0.345187 0.21 0.381937 0.231 ;
  RECT 0.381937 0.191625 0.549935 0.21 ;
      LAYER M1 ;
  RECT 0.0538125 0.418687 0.179812 0.437063 ;
  RECT 0.179812 0.108937 0.242812 0.127312 ;
  RECT 0.179812 0.418687 0.242812 0.437063 ;
  RECT 0.242812 0.108937 0.261188 0.127312 ;
  RECT 0.242812 0.127312 0.261188 0.254625 ;
  RECT 0.242812 0.254625 0.261188 0.271688 ;
  RECT 0.242812 0.271688 0.261188 0.300563 ;
  RECT 0.242812 0.300563 0.261188 0.418687 ;
  RECT 0.242812 0.418687 0.261188 0.437063 ;
  RECT 0.261188 0.418687 0.345187 0.437063 ;
  RECT 0.345187 0.254625 0.381937 0.271688 ;
  RECT 0.345187 0.271688 0.381937 0.300563 ;
  RECT 0.345187 0.300563 0.381937 0.418687 ;
  RECT 0.345187 0.418687 0.381937 0.437063 ;
  RECT 0.381937 0.271688 0.53412 0.300563 ;
  RECT 0.0328125 0.063 0.0511875 0.20475 ;
  RECT 0.0328125 0.20475 0.0511875 0.223125 ;
  RECT 0.0328125 0.223125 0.0511875 0.265125 ;
  RECT 0.0328125 0.265125 0.0511875 0.389813 ;
  RECT 0.0511875 0.20475 0.116812 0.223125 ;
  RECT 0.116812 0.20475 0.135187 0.223125 ;
  RECT 0.116812 0.223125 0.135187 0.265125 ;
  RECT 0.0958125 0.372685 0.132562 0.395062 ;
  RECT 0.132562 0.066872 0.150937 0.0853125 ;
  RECT 0.132562 0.0853125 0.150937 0.150937 ;
  RECT 0.132562 0.150937 0.150937 0.169312 ;
  RECT 0.132562 0.372685 0.150937 0.395062 ;
  RECT 0.150937 0.066872 0.200812 0.0853125 ;
  RECT 0.150937 0.150937 0.200812 0.169312 ;
  RECT 0.150937 0.372685 0.200812 0.395062 ;
  RECT 0.200812 0.066872 0.219187 0.0853125 ;
  RECT 0.200812 0.150937 0.219187 0.169312 ;
  RECT 0.200812 0.169312 0.219187 0.191625 ;
  RECT 0.200812 0.191625 0.219187 0.21 ;
  RECT 0.200812 0.21 0.219187 0.231 ;
  RECT 0.200812 0.231 0.219187 0.372685 ;
  RECT 0.200812 0.372685 0.219187 0.395062 ;
  RECT 0.219187 0.066872 0.345187 0.0853125 ;
  RECT 0.345187 0.066872 0.381937 0.0853125 ;
  RECT 0.345187 0.0853125 0.381937 0.150937 ;
  RECT 0.345187 0.150937 0.381937 0.169312 ;
  RECT 0.345187 0.169312 0.381937 0.191625 ;
  RECT 0.345187 0.191625 0.381937 0.21 ;
  RECT 0.345187 0.21 0.381937 0.231 ;
  RECT 0.381937 0.191625 0.549935 0.21 ;
  END
END TBUF_X4

MACRO TBUF_X8
  CLASS core ;
  FOREIGN TBUF_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.882 BY 0.504 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.252 0.093122 0.317625 ;
  RECT 0.0748125 0.317625 0.093122 0.336 ;
  RECT 0.093122 0.317625 0.145687 0.336 ;
  RECT 0.145687 0.317625 0.200812 0.336 ;
  RECT 0.200812 0.21 0.219187 0.252 ;
  RECT 0.200812 0.252 0.219187 0.317625 ;
  RECT 0.200812 0.317625 0.219187 0.336 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.326813 0.226997 0.345187 0.263813 ;
  RECT 0.326813 0.263813 0.345187 0.284813 ;
  RECT 0.326813 0.284813 0.345187 0.378 ;
  RECT 0.345187 0.263813 0.408187 0.284813 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.535435 0.042 0.5565 0.0872815 ;
  RECT 0.535435 0.0872815 0.5565 0.105 ;
  RECT 0.535435 0.105 0.5565 0.126 ;
  RECT 0.535435 0.340595 0.5565 0.378655 ;
  RECT 0.535435 0.378655 0.5565 0.379312 ;
  RECT 0.535435 0.379312 0.5565 0.462 ;
  RECT 0.5565 0.105 0.776345 0.126 ;
  RECT 0.5565 0.340595 0.776345 0.378655 ;
  RECT 0.776345 0.105 0.78619 0.126 ;
  RECT 0.776345 0.340595 0.78619 0.378655 ;
  RECT 0.78619 0.105 0.7875 0.126 ;
  RECT 0.78619 0.340595 0.7875 0.378655 ;
  RECT 0.7875 0.042 0.8085 0.0872815 ;
  RECT 0.7875 0.0872815 0.8085 0.105 ;
  RECT 0.7875 0.105 0.8085 0.126 ;
  RECT 0.7875 0.340595 0.8085 0.378655 ;
  RECT 0.7875 0.378655 0.8085 0.379312 ;
  RECT 0.7875 0.379312 0.8085 0.462 ;
  RECT 0.8085 0.0872815 0.83081 0.105 ;
  RECT 0.8085 0.105 0.83081 0.126 ;
  RECT 0.8085 0.340595 0.83081 0.378655 ;
  RECT 0.8085 0.378655 0.83081 0.379312 ;
  RECT 0.83081 0.0872815 0.849185 0.105 ;
  RECT 0.83081 0.105 0.849185 0.126 ;
  RECT 0.83081 0.126 0.849185 0.340595 ;
  RECT 0.83081 0.340595 0.849185 0.378655 ;
  RECT 0.83081 0.378655 0.849185 0.379312 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.776345 0.522375 ;
  RECT 0.776345 0.485625 0.78619 0.522375 ;
  RECT 0.78619 0.485625 0.888565 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.888565 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0328125 0.04725 0.0511875 0.20475 ;
  RECT 0.0328125 0.20475 0.0511875 0.223125 ;
  RECT 0.0328125 0.223125 0.0511875 0.282187 ;
  RECT 0.0328125 0.282187 0.0511875 0.418687 ;
  RECT 0.0511875 0.20475 0.116812 0.223125 ;
  RECT 0.116812 0.20475 0.145687 0.223125 ;
  RECT 0.116812 0.223125 0.145687 0.282187 ;
  RECT 0.0958125 0.376688 0.132562 0.395062 ;
  RECT 0.132562 0.066872 0.150937 0.0853125 ;
  RECT 0.132562 0.0853125 0.150937 0.150937 ;
  RECT 0.132562 0.150937 0.150937 0.169312 ;
  RECT 0.132562 0.376688 0.150937 0.395062 ;
  RECT 0.150937 0.066872 0.242812 0.0853125 ;
  RECT 0.150937 0.150937 0.242812 0.169312 ;
  RECT 0.150937 0.376688 0.242812 0.395062 ;
  RECT 0.242812 0.066872 0.261188 0.0853125 ;
  RECT 0.242812 0.150937 0.261188 0.169312 ;
  RECT 0.242812 0.169312 0.261188 0.187622 ;
  RECT 0.242812 0.187622 0.261188 0.224437 ;
  RECT 0.242812 0.224437 0.261188 0.376688 ;
  RECT 0.242812 0.376688 0.261188 0.395062 ;
  RECT 0.261188 0.066872 0.452748 0.0853125 ;
  RECT 0.452748 0.066872 0.471187 0.0853125 ;
  RECT 0.452748 0.0853125 0.471187 0.150937 ;
  RECT 0.452748 0.150937 0.471187 0.169312 ;
  RECT 0.452748 0.169312 0.471187 0.187622 ;
  RECT 0.452748 0.187622 0.471187 0.224437 ;
  RECT 0.471187 0.169312 0.78619 0.187622 ;
  RECT 0.0800625 0.418687 0.179812 0.437063 ;
  RECT 0.179812 0.108937 0.284813 0.127312 ;
  RECT 0.179812 0.418687 0.284813 0.437063 ;
  RECT 0.284813 0.108937 0.303187 0.127312 ;
  RECT 0.284813 0.127312 0.303187 0.253312 ;
  RECT 0.284813 0.253312 0.303187 0.26447 ;
  RECT 0.284813 0.26447 0.303187 0.30253 ;
  RECT 0.284813 0.30253 0.303187 0.418687 ;
  RECT 0.284813 0.418687 0.303187 0.437063 ;
  RECT 0.303187 0.418687 0.433125 0.437063 ;
  RECT 0.433125 0.253312 0.471187 0.26447 ;
  RECT 0.433125 0.26447 0.471187 0.30253 ;
  RECT 0.433125 0.30253 0.471187 0.418687 ;
  RECT 0.433125 0.418687 0.471187 0.437063 ;
  RECT 0.471187 0.26447 0.776345 0.30253 ;
      LAYER M1 ;
  RECT 0.0328125 0.04725 0.0511875 0.20475 ;
  RECT 0.0328125 0.20475 0.0511875 0.223125 ;
  RECT 0.0328125 0.223125 0.0511875 0.282187 ;
  RECT 0.0328125 0.282187 0.0511875 0.418687 ;
  RECT 0.0511875 0.20475 0.116812 0.223125 ;
  RECT 0.116812 0.20475 0.145687 0.223125 ;
  RECT 0.116812 0.223125 0.145687 0.282187 ;
  RECT 0.0958125 0.376688 0.132562 0.395062 ;
  RECT 0.132562 0.066872 0.150937 0.0853125 ;
  RECT 0.132562 0.0853125 0.150937 0.150937 ;
  RECT 0.132562 0.150937 0.150937 0.169312 ;
  RECT 0.132562 0.376688 0.150937 0.395062 ;
  RECT 0.150937 0.066872 0.242812 0.0853125 ;
  RECT 0.150937 0.150937 0.242812 0.169312 ;
  RECT 0.150937 0.376688 0.242812 0.395062 ;
  RECT 0.242812 0.066872 0.261188 0.0853125 ;
  RECT 0.242812 0.150937 0.261188 0.169312 ;
  RECT 0.242812 0.169312 0.261188 0.187622 ;
  RECT 0.242812 0.187622 0.261188 0.224437 ;
  RECT 0.242812 0.224437 0.261188 0.376688 ;
  RECT 0.242812 0.376688 0.261188 0.395062 ;
  RECT 0.261188 0.066872 0.452748 0.0853125 ;
  RECT 0.452748 0.066872 0.471187 0.0853125 ;
  RECT 0.452748 0.0853125 0.471187 0.150937 ;
  RECT 0.452748 0.150937 0.471187 0.169312 ;
  RECT 0.452748 0.169312 0.471187 0.187622 ;
  RECT 0.452748 0.187622 0.471187 0.224437 ;
  RECT 0.471187 0.169312 0.78619 0.187622 ;
  RECT 0.0800625 0.418687 0.179812 0.437063 ;
  RECT 0.179812 0.108937 0.284813 0.127312 ;
  RECT 0.179812 0.418687 0.284813 0.437063 ;
  RECT 0.284813 0.108937 0.303187 0.127312 ;
  RECT 0.284813 0.127312 0.303187 0.253312 ;
  RECT 0.284813 0.253312 0.303187 0.26447 ;
  RECT 0.284813 0.26447 0.303187 0.30253 ;
  RECT 0.284813 0.30253 0.303187 0.418687 ;
  RECT 0.284813 0.418687 0.303187 0.437063 ;
  RECT 0.303187 0.418687 0.433125 0.437063 ;
  RECT 0.433125 0.253312 0.471187 0.26447 ;
  RECT 0.433125 0.26447 0.471187 0.30253 ;
  RECT 0.433125 0.30253 0.471187 0.418687 ;
  RECT 0.433125 0.418687 0.471187 0.437063 ;
  RECT 0.471187 0.26447 0.776345 0.30253 ;
  END
END TBUF_X8

MACRO TBUF_X12
  CLASS core ;
  FOREIGN TBUF_X12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 1.134 BY 0.504 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.252 0.093122 0.334688 ;
  RECT 0.0748125 0.334688 0.093122 0.353063 ;
  RECT 0.093122 0.334688 0.135187 0.353063 ;
  RECT 0.135187 0.334688 0.158812 0.353063 ;
  RECT 0.158812 0.200812 0.177187 0.252 ;
  RECT 0.158812 0.252 0.177187 0.334688 ;
  RECT 0.158812 0.334688 0.177187 0.353063 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.284813 0.263813 0.326813 0.294 ;
  RECT 0.326813 0.226997 0.345187 0.263813 ;
  RECT 0.326813 0.263813 0.345187 0.294 ;
  RECT 0.345187 0.263813 0.410813 0.294 ;
  RECT 0.410813 0.263813 0.429187 0.294 ;
  RECT 0.410813 0.294 0.429187 0.378 ;
  RECT 0.429187 0.263813 0.465938 0.294 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 1.10512 0.522375 ;
  RECT 1.10512 0.485625 1.14056 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 1.14056 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0958125 0.418687 0.179812 0.437063 ;
  RECT 0.179812 0.108937 0.242812 0.127312 ;
  RECT 0.179812 0.418687 0.242812 0.437063 ;
  RECT 0.242812 0.108937 0.261188 0.127312 ;
  RECT 0.242812 0.127312 0.261188 0.233625 ;
  RECT 0.242812 0.233625 0.261188 0.248062 ;
  RECT 0.242812 0.248062 0.261188 0.279562 ;
  RECT 0.242812 0.279562 0.261188 0.418687 ;
  RECT 0.242812 0.418687 0.261188 0.437063 ;
  RECT 0.261188 0.418687 0.513845 0.437063 ;
  RECT 0.513845 0.233625 0.550595 0.248062 ;
  RECT 0.513845 0.248062 0.550595 0.279562 ;
  RECT 0.513845 0.279562 0.550595 0.418687 ;
  RECT 0.513845 0.418687 0.550595 0.437063 ;
  RECT 0.550595 0.248062 1.02178 0.279562 ;
  RECT 0.57881 0.066872 0.61097 0.0853125 ;
  RECT 0.61097 0.066872 0.64903 0.0853125 ;
  RECT 0.61097 0.349125 0.64903 0.37006 ;
  RECT 0.61097 0.37006 0.64903 0.406875 ;
  RECT 0.64903 0.066872 1.03162 0.0853125 ;
  RECT 0.64903 0.349125 1.03162 0.37006 ;
  RECT 1.03162 0.0479062 1.04081 0.066872 ;
  RECT 1.03162 0.066872 1.04081 0.0853125 ;
  RECT 1.03162 0.349125 1.04081 0.37006 ;
  RECT 1.04081 0.0479062 1.05919 0.066872 ;
  RECT 1.04081 0.066872 1.05919 0.0853125 ;
  RECT 1.04081 0.349125 1.05919 0.37006 ;
  RECT 1.04081 0.37006 1.05919 0.406875 ;
  RECT 1.04081 0.406875 1.05919 0.4095 ;
  RECT 1.05919 0.0479062 1.06831 0.066872 ;
  RECT 1.05919 0.066872 1.06831 0.0853125 ;
  RECT 1.05919 0.349125 1.06831 0.37006 ;
  RECT 1.06831 0.066872 1.06903 0.0853125 ;
  RECT 1.06831 0.349125 1.06903 0.37006 ;
  RECT 1.06903 0.066872 1.10512 0.0853125 ;
  RECT 1.06903 0.0853125 1.10512 0.349125 ;
  RECT 1.06903 0.349125 1.10512 0.37006 ;
  RECT 0.0328125 0.114122 0.0511875 0.20475 ;
  RECT 0.0328125 0.20475 0.0511875 0.223125 ;
  RECT 0.0328125 0.223125 0.0511875 0.265125 ;
  RECT 0.0328125 0.265125 0.0511875 0.441 ;
  RECT 0.0511875 0.20475 0.116812 0.223125 ;
  RECT 0.116812 0.20475 0.135187 0.223125 ;
  RECT 0.116812 0.223125 0.135187 0.265125 ;
  RECT 0.093122 0.066872 0.0958125 0.0853125 ;
  RECT 0.093122 0.0853125 0.0958125 0.150937 ;
  RECT 0.093122 0.150937 0.0958125 0.164062 ;
  RECT 0.093122 0.164062 0.0958125 0.169312 ;
  RECT 0.0958125 0.066872 0.111562 0.0853125 ;
  RECT 0.0958125 0.0853125 0.111562 0.150937 ;
  RECT 0.0958125 0.150937 0.111562 0.164062 ;
  RECT 0.0958125 0.164062 0.111562 0.169312 ;
  RECT 0.0958125 0.376688 0.111562 0.395062 ;
  RECT 0.111562 0.066872 0.200812 0.0853125 ;
  RECT 0.111562 0.150937 0.200812 0.164062 ;
  RECT 0.111562 0.164062 0.200812 0.169312 ;
  RECT 0.111562 0.376688 0.200812 0.395062 ;
  RECT 0.200812 0.066872 0.219187 0.0853125 ;
  RECT 0.200812 0.150937 0.219187 0.164062 ;
  RECT 0.200812 0.164062 0.219187 0.169312 ;
  RECT 0.200812 0.169312 0.219187 0.192937 ;
  RECT 0.200812 0.192937 0.219187 0.376688 ;
  RECT 0.200812 0.376688 0.219187 0.395062 ;
  RECT 0.219187 0.066872 0.51319 0.0853125 ;
  RECT 0.51319 0.066872 0.53412 0.0853125 ;
  RECT 0.51319 0.0853125 0.53412 0.150937 ;
  RECT 0.51319 0.150937 0.53412 0.164062 ;
  RECT 0.51319 0.164062 0.53412 0.169312 ;
  RECT 0.51319 0.169312 0.53412 0.192937 ;
  RECT 0.53412 0.164062 1.04541 0.169312 ;
  RECT 0.53412 0.169312 1.04541 0.192937 ;
      LAYER M1 ;
  RECT 0.0958125 0.418687 0.179812 0.437063 ;
  RECT 0.179812 0.108937 0.242812 0.127312 ;
  RECT 0.179812 0.418687 0.242812 0.437063 ;
  RECT 0.242812 0.108937 0.261188 0.127312 ;
  RECT 0.242812 0.127312 0.261188 0.233625 ;
  RECT 0.242812 0.233625 0.261188 0.248062 ;
  RECT 0.242812 0.248062 0.261188 0.279562 ;
  RECT 0.242812 0.279562 0.261188 0.418687 ;
  RECT 0.242812 0.418687 0.261188 0.437063 ;
  RECT 0.261188 0.418687 0.513845 0.437063 ;
  RECT 0.513845 0.233625 0.550595 0.248062 ;
  RECT 0.513845 0.248062 0.550595 0.279562 ;
  RECT 0.513845 0.279562 0.550595 0.418687 ;
  RECT 0.513845 0.418687 0.550595 0.437063 ;
  RECT 0.550595 0.248062 1.02178 0.279562 ;
  RECT 0.57881 0.066872 0.61097 0.0853125 ;
  RECT 0.61097 0.066872 0.64903 0.0853125 ;
  RECT 0.61097 0.349125 0.64903 0.37006 ;
  RECT 0.61097 0.37006 0.64903 0.406875 ;
  RECT 0.64903 0.066872 1.03162 0.0853125 ;
  RECT 0.64903 0.349125 1.03162 0.37006 ;
  RECT 1.03162 0.0479062 1.04081 0.066872 ;
  RECT 1.03162 0.066872 1.04081 0.0853125 ;
  RECT 1.03162 0.349125 1.04081 0.37006 ;
  RECT 1.04081 0.0479062 1.05919 0.066872 ;
  RECT 1.04081 0.066872 1.05919 0.0853125 ;
  RECT 1.04081 0.349125 1.05919 0.37006 ;
  RECT 1.04081 0.37006 1.05919 0.406875 ;
  RECT 1.04081 0.406875 1.05919 0.4095 ;
  RECT 1.05919 0.0479062 1.06831 0.066872 ;
  RECT 1.05919 0.066872 1.06831 0.0853125 ;
  RECT 1.05919 0.349125 1.06831 0.37006 ;
  RECT 1.06831 0.066872 1.06903 0.0853125 ;
  RECT 1.06831 0.349125 1.06903 0.37006 ;
  RECT 1.06903 0.066872 1.10512 0.0853125 ;
  RECT 1.06903 0.0853125 1.10512 0.349125 ;
  RECT 1.06903 0.349125 1.10512 0.37006 ;
  RECT 0.0328125 0.114122 0.0511875 0.20475 ;
  RECT 0.0328125 0.20475 0.0511875 0.223125 ;
  RECT 0.0328125 0.223125 0.0511875 0.265125 ;
  RECT 0.0328125 0.265125 0.0511875 0.441 ;
  RECT 0.0511875 0.20475 0.116812 0.223125 ;
  RECT 0.116812 0.20475 0.135187 0.223125 ;
  RECT 0.116812 0.223125 0.135187 0.265125 ;
  RECT 0.093122 0.066872 0.0958125 0.0853125 ;
  RECT 0.093122 0.0853125 0.0958125 0.150937 ;
  RECT 0.093122 0.150937 0.0958125 0.164062 ;
  RECT 0.093122 0.164062 0.0958125 0.169312 ;
  RECT 0.0958125 0.066872 0.111562 0.0853125 ;
  RECT 0.0958125 0.0853125 0.111562 0.150937 ;
  RECT 0.0958125 0.150937 0.111562 0.164062 ;
  RECT 0.0958125 0.164062 0.111562 0.169312 ;
  RECT 0.0958125 0.376688 0.111562 0.395062 ;
  RECT 0.111562 0.066872 0.200812 0.0853125 ;
  RECT 0.111562 0.150937 0.200812 0.164062 ;
  RECT 0.111562 0.164062 0.200812 0.169312 ;
  RECT 0.111562 0.376688 0.200812 0.395062 ;
  RECT 0.200812 0.066872 0.219187 0.0853125 ;
  RECT 0.200812 0.150937 0.219187 0.164062 ;
  RECT 0.200812 0.164062 0.219187 0.169312 ;
  RECT 0.200812 0.169312 0.219187 0.192937 ;
  RECT 0.200812 0.192937 0.219187 0.376688 ;
  RECT 0.200812 0.376688 0.219187 0.395062 ;
  RECT 0.219187 0.066872 0.51319 0.0853125 ;
  RECT 0.51319 0.066872 0.53412 0.0853125 ;
  RECT 0.51319 0.0853125 0.53412 0.150937 ;
  RECT 0.51319 0.150937 0.53412 0.164062 ;
  RECT 0.51319 0.164062 0.53412 0.169312 ;
  RECT 0.51319 0.169312 0.53412 0.192937 ;
  RECT 0.53412 0.164062 1.04541 0.169312 ;
  RECT 0.53412 0.169312 1.04541 0.192937 ;
  END
END TBUF_X12

MACRO TBUF_X16
  CLASS core ;
  FOREIGN TBUF_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 1.386 BY 0.504 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0748125 0.255937 0.093122 0.318937 ;
  RECT 0.0748125 0.318937 0.093122 0.337313 ;
  RECT 0.093122 0.318937 0.114122 0.337313 ;
  RECT 0.114122 0.318937 0.1575 0.337313 ;
  RECT 0.1575 0.21 0.1785 0.255937 ;
  RECT 0.1575 0.255937 0.1785 0.318937 ;
  RECT 0.1575 0.318937 0.1785 0.337313 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.303187 0.263813 0.368812 0.294 ;
  RECT 0.368812 0.226997 0.387188 0.263813 ;
  RECT 0.368812 0.263813 0.387188 0.294 ;
  RECT 0.387188 0.263813 0.452748 0.294 ;
  RECT 0.452748 0.263813 0.471187 0.294 ;
  RECT 0.452748 0.294 0.471187 0.378 ;
  RECT 0.471187 0.263813 0.59194 0.294 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.7035 0.042 0.7245 0.093122 ;
  RECT 0.7035 0.093122 0.7245 0.13125 ;
  RECT 0.7035 0.34125 0.7245 0.378 ;
  RECT 0.7035 0.378 0.7245 0.462 ;
  RECT 0.7245 0.093122 1.2915 0.13125 ;
  RECT 0.7245 0.34125 1.2915 0.378 ;
  RECT 1.2915 0.042 1.29937 0.093122 ;
  RECT 1.2915 0.093122 1.29937 0.13125 ;
  RECT 1.2915 0.34125 1.29937 0.378 ;
  RECT 1.2915 0.378 1.29937 0.462 ;
  RECT 1.29937 0.042 1.31119 0.093122 ;
  RECT 1.29937 0.093122 1.31119 0.13125 ;
  RECT 1.29937 0.34125 1.31119 0.378 ;
  RECT 1.29937 0.378 1.31119 0.462 ;
  RECT 1.31119 0.042 1.3125 0.093122 ;
  RECT 1.31119 0.093122 1.3125 0.13125 ;
  RECT 1.31119 0.34125 1.3125 0.378 ;
  RECT 1.31119 0.378 1.3125 0.462 ;
  RECT 1.3125 0.093122 1.33475 0.13125 ;
  RECT 1.3125 0.34125 1.33475 0.378 ;
  RECT 1.33475 0.093122 1.35319 0.13125 ;
  RECT 1.33475 0.13125 1.35319 0.34125 ;
  RECT 1.33475 0.34125 1.35319 0.378 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 1.29937 0.522375 ;
  RECT 1.29937 0.485625 1.31119 0.522375 ;
  RECT 1.31119 0.485625 1.39256 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 1.39256 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0328125 0.04725 0.0511875 0.171937 ;
  RECT 0.0328125 0.171937 0.0511875 0.190312 ;
  RECT 0.0328125 0.190312 0.0511875 0.226997 ;
  RECT 0.0328125 0.226997 0.0511875 0.39375 ;
  RECT 0.0511875 0.171937 0.093122 0.190312 ;
  RECT 0.093122 0.171937 0.114122 0.190312 ;
  RECT 0.093122 0.190312 0.114122 0.226997 ;
  RECT 0.0958125 0.418687 0.179812 0.437063 ;
  RECT 0.179812 0.108937 0.261188 0.129937 ;
  RECT 0.179812 0.418687 0.261188 0.437063 ;
  RECT 0.261188 0.108937 0.279562 0.129937 ;
  RECT 0.261188 0.129937 0.279562 0.26447 ;
  RECT 0.261188 0.26447 0.279562 0.30253 ;
  RECT 0.261188 0.30253 0.279562 0.418687 ;
  RECT 0.261188 0.418687 0.279562 0.437063 ;
  RECT 0.279562 0.418687 0.62081 0.437063 ;
  RECT 0.62081 0.26447 0.63919 0.30253 ;
  RECT 0.62081 0.30253 0.63919 0.418687 ;
  RECT 0.62081 0.418687 0.63919 0.437063 ;
  RECT 0.63919 0.26447 1.29937 0.30253 ;
  RECT 0.0958125 0.372685 0.137812 0.395062 ;
  RECT 0.137812 0.066872 0.156187 0.0853125 ;
  RECT 0.137812 0.0853125 0.156187 0.153562 ;
  RECT 0.137812 0.153562 0.156187 0.171937 ;
  RECT 0.137812 0.372685 0.156187 0.395062 ;
  RECT 0.156187 0.066872 0.213937 0.0853125 ;
  RECT 0.156187 0.153562 0.213937 0.171937 ;
  RECT 0.156187 0.372685 0.213937 0.395062 ;
  RECT 0.213937 0.066872 0.237562 0.0853125 ;
  RECT 0.213937 0.153562 0.237562 0.171937 ;
  RECT 0.213937 0.171937 0.237562 0.179156 ;
  RECT 0.213937 0.179156 0.237562 0.217219 ;
  RECT 0.213937 0.217219 0.237562 0.372685 ;
  RECT 0.213937 0.372685 0.237562 0.395062 ;
  RECT 0.237562 0.066872 0.62081 0.0853125 ;
  RECT 0.62081 0.066872 0.63919 0.0853125 ;
  RECT 0.62081 0.0853125 0.63919 0.153562 ;
  RECT 0.62081 0.153562 0.63919 0.171937 ;
  RECT 0.62081 0.171937 0.63919 0.179156 ;
  RECT 0.62081 0.179156 0.63919 0.217219 ;
  RECT 0.63919 0.179156 1.31119 0.217219 ;
      LAYER M1 ;
  RECT 0.0328125 0.04725 0.0511875 0.171937 ;
  RECT 0.0328125 0.171937 0.0511875 0.190312 ;
  RECT 0.0328125 0.190312 0.0511875 0.226997 ;
  RECT 0.0328125 0.226997 0.0511875 0.39375 ;
  RECT 0.0511875 0.171937 0.093122 0.190312 ;
  RECT 0.093122 0.171937 0.114122 0.190312 ;
  RECT 0.093122 0.190312 0.114122 0.226997 ;
  RECT 0.0958125 0.418687 0.179812 0.437063 ;
  RECT 0.179812 0.108937 0.261188 0.129937 ;
  RECT 0.179812 0.418687 0.261188 0.437063 ;
  RECT 0.261188 0.108937 0.279562 0.129937 ;
  RECT 0.261188 0.129937 0.279562 0.26447 ;
  RECT 0.261188 0.26447 0.279562 0.30253 ;
  RECT 0.261188 0.30253 0.279562 0.418687 ;
  RECT 0.261188 0.418687 0.279562 0.437063 ;
  RECT 0.279562 0.418687 0.62081 0.437063 ;
  RECT 0.62081 0.26447 0.63919 0.30253 ;
  RECT 0.62081 0.30253 0.63919 0.418687 ;
  RECT 0.62081 0.418687 0.63919 0.437063 ;
  RECT 0.63919 0.26447 1.29937 0.30253 ;
  RECT 0.0958125 0.372685 0.137812 0.395062 ;
  RECT 0.137812 0.066872 0.156187 0.0853125 ;
  RECT 0.137812 0.0853125 0.156187 0.153562 ;
  RECT 0.137812 0.153562 0.156187 0.171937 ;
  RECT 0.137812 0.372685 0.156187 0.395062 ;
  RECT 0.156187 0.066872 0.213937 0.0853125 ;
  RECT 0.156187 0.153562 0.213937 0.171937 ;
  RECT 0.156187 0.372685 0.213937 0.395062 ;
  RECT 0.213937 0.066872 0.237562 0.0853125 ;
  RECT 0.213937 0.153562 0.237562 0.171937 ;
  RECT 0.213937 0.171937 0.237562 0.179156 ;
  RECT 0.213937 0.179156 0.237562 0.217219 ;
  RECT 0.213937 0.217219 0.237562 0.372685 ;
  RECT 0.213937 0.372685 0.237562 0.395062 ;
  RECT 0.237562 0.066872 0.62081 0.0853125 ;
  RECT 0.62081 0.066872 0.63919 0.0853125 ;
  RECT 0.62081 0.0853125 0.63919 0.153562 ;
  RECT 0.62081 0.153562 0.63919 0.171937 ;
  RECT 0.62081 0.171937 0.63919 0.179156 ;
  RECT 0.62081 0.179156 0.63919 0.217219 ;
  RECT 0.63919 0.179156 1.31119 0.217219 ;
  END
END TBUF_X16

MACRO TIEH
  CLASS core ;
  FOREIGN TIEH 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.126 BY 0.504 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0715315 0.310405 0.093122 0.462 ;
  RECT 0.093122 0.310405 0.096469 0.462 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.093122 0.522375 ;
  RECT 0.093122 0.485625 0.132562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.132562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0748125 0.063 0.093122 0.28153 ;
      LAYER M1 ;
  RECT 0.0748125 0.063 0.093122 0.28153 ;
  END
END TIEH

MACRO TIEL
  CLASS core ;
  FOREIGN TIEL 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.126 BY 0.504 ;
  PIN Z
    DIRECTION INOUT ;
    PORT
      LAYER M1 ;
  RECT 0.0715315 0.042 0.096469 0.174562 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.093122 0.522375 ;
  RECT 0.093122 0.485625 0.132562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.132562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.0748125 0.2205 0.093122 0.441 ;
      LAYER M1 ;
  RECT 0.0748125 0.2205 0.093122 0.441 ;
  END
END TIEL

MACRO XNOR2_X1
  CLASS core ;
  FOREIGN XNOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.378 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.165375 0.137812 0.18375 ;
  RECT 0.116812 0.18375 0.137812 0.280875 ;
  RECT 0.137812 0.165375 0.242812 0.18375 ;
  RECT 0.242812 0.165375 0.261188 0.18375 ;
  RECT 0.242812 0.18375 0.261188 0.280875 ;
  RECT 0.242812 0.280875 0.261188 0.294 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.158812 0.0511875 0.21 ;
  RECT 0.0328125 0.21 0.0511875 0.443625 ;
  RECT 0.0328125 0.443625 0.0511875 0.462 ;
  RECT 0.0511875 0.443625 0.179812 0.462 ;
  RECT 0.179812 0.443625 0.326813 0.462 ;
  RECT 0.326813 0.21 0.345187 0.443625 ;
  RECT 0.326813 0.443625 0.345187 0.462 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.182437 0.358312 0.198187 0.35897 ;
  RECT 0.182437 0.35897 0.198187 0.394405 ;
  RECT 0.182437 0.394405 0.198187 0.395062 ;
  RECT 0.198187 0.108937 0.219187 0.127312 ;
  RECT 0.198187 0.358312 0.219187 0.35897 ;
  RECT 0.198187 0.35897 0.219187 0.394405 ;
  RECT 0.198187 0.394405 0.219187 0.395062 ;
  RECT 0.219187 0.108937 0.284813 0.127312 ;
  RECT 0.219187 0.35897 0.284813 0.394405 ;
  RECT 0.284813 0.108937 0.303187 0.127312 ;
  RECT 0.284813 0.16275 0.303187 0.181125 ;
  RECT 0.284813 0.181125 0.303187 0.358312 ;
  RECT 0.284813 0.358312 0.303187 0.35897 ;
  RECT 0.284813 0.35897 0.303187 0.394405 ;
  RECT 0.303187 0.108937 0.32353 0.127312 ;
  RECT 0.303187 0.16275 0.32353 0.181125 ;
  RECT 0.32353 0.108937 0.34847 0.127312 ;
  RECT 0.32353 0.127312 0.34847 0.16275 ;
  RECT 0.32353 0.16275 0.34847 0.181125 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.179812 0.522375 ;
  RECT 0.179812 0.485625 0.351095 0.522375 ;
  RECT 0.351095 0.485625 0.384562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.384562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.137812 0.066872 0.351095 0.0853125 ;
  RECT 0.0748125 0.12075 0.093122 0.14175 ;
  RECT 0.0748125 0.14175 0.093122 0.223125 ;
  RECT 0.0748125 0.223125 0.093122 0.3045 ;
  RECT 0.0748125 0.3045 0.093122 0.322875 ;
  RECT 0.0748125 0.322875 0.093122 0.36225 ;
  RECT 0.093122 0.12075 0.153562 0.14175 ;
  RECT 0.093122 0.3045 0.153562 0.322875 ;
  RECT 0.153562 0.3045 0.161437 0.322875 ;
  RECT 0.161437 0.223125 0.179812 0.3045 ;
  RECT 0.161437 0.3045 0.179812 0.322875 ;
      LAYER M1 ;
  RECT 0.137812 0.066872 0.351095 0.0853125 ;
  RECT 0.0748125 0.12075 0.093122 0.14175 ;
  RECT 0.0748125 0.14175 0.093122 0.223125 ;
  RECT 0.0748125 0.223125 0.093122 0.3045 ;
  RECT 0.0748125 0.3045 0.093122 0.322875 ;
  RECT 0.0748125 0.322875 0.093122 0.36225 ;
  RECT 0.093122 0.12075 0.153562 0.14175 ;
  RECT 0.093122 0.3045 0.153562 0.322875 ;
  RECT 0.153562 0.3045 0.161437 0.322875 ;
  RECT 0.161437 0.223125 0.179812 0.3045 ;
  RECT 0.161437 0.3045 0.179812 0.322875 ;
  END
END XNOR2_X1

MACRO XOR2_X1
  CLASS core ;
  FOREIGN XOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CORE_TypTyp_0p4_25 ;
SIZE 0.378 BY 0.504 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.116812 0.225684 0.137812 0.318937 ;
  RECT 0.116812 0.318937 0.137812 0.337313 ;
  RECT 0.137812 0.318937 0.179812 0.337313 ;
  RECT 0.179812 0.318937 0.242812 0.337313 ;
  RECT 0.242812 0.21 0.261188 0.225684 ;
  RECT 0.242812 0.225684 0.261188 0.318937 ;
  RECT 0.242812 0.318937 0.261188 0.337313 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
  RECT 0.0328125 0.042 0.0511875 0.060375 ;
  RECT 0.0328125 0.060375 0.0511875 0.294 ;
  RECT 0.0328125 0.294 0.0511875 0.345187 ;
  RECT 0.0511875 0.042 0.326813 0.060375 ;
  RECT 0.326813 0.042 0.345187 0.060375 ;
  RECT 0.326813 0.060375 0.345187 0.294 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
  RECT 0.180469 0.106969 0.206719 0.107625 ;
  RECT 0.180469 0.107625 0.206719 0.145687 ;
  RECT 0.206719 0.106969 0.219187 0.107625 ;
  RECT 0.206719 0.107625 0.219187 0.145687 ;
  RECT 0.206719 0.376688 0.219187 0.395062 ;
  RECT 0.219187 0.107625 0.284813 0.145687 ;
  RECT 0.219187 0.376688 0.284813 0.395062 ;
  RECT 0.284813 0.107625 0.303187 0.145687 ;
  RECT 0.284813 0.145687 0.303187 0.322875 ;
  RECT 0.284813 0.322875 0.303187 0.34125 ;
  RECT 0.284813 0.376688 0.303187 0.395062 ;
  RECT 0.303187 0.322875 0.3255 0.34125 ;
  RECT 0.303187 0.376688 0.3255 0.395062 ;
  RECT 0.3255 0.322875 0.3465 0.34125 ;
  RECT 0.3255 0.34125 0.3465 0.376688 ;
  RECT 0.3255 0.376688 0.3465 0.395062 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 0.485625 0.351095 0.522375 ;
  RECT 0.351095 0.485625 0.384562 0.522375 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
  RECT -0.0065625 -0.018375 0.384562 0.018375 ;
    END
  END VSS
  OBS
      LAYER M1 ;
  RECT 0.161437 0.418687 0.351095 0.437063 ;
  RECT 0.0748125 0.08925 0.093122 0.18375 ;
  RECT 0.0748125 0.18375 0.093122 0.202125 ;
  RECT 0.0748125 0.202125 0.093122 0.2835 ;
  RECT 0.0748125 0.2835 0.093122 0.36225 ;
  RECT 0.0748125 0.36225 0.093122 0.38325 ;
  RECT 0.093122 0.18375 0.161437 0.202125 ;
  RECT 0.093122 0.36225 0.161437 0.38325 ;
  RECT 0.161437 0.18375 0.162094 0.202125 ;
  RECT 0.161437 0.202125 0.162094 0.2835 ;
  RECT 0.161437 0.36225 0.162094 0.38325 ;
  RECT 0.162094 0.18375 0.179812 0.202125 ;
  RECT 0.162094 0.202125 0.179812 0.2835 ;
      LAYER M1 ;
  RECT 0.161437 0.418687 0.351095 0.437063 ;
  RECT 0.0748125 0.08925 0.093122 0.18375 ;
  RECT 0.0748125 0.18375 0.093122 0.202125 ;
  RECT 0.0748125 0.202125 0.093122 0.2835 ;
  RECT 0.0748125 0.2835 0.093122 0.36225 ;
  RECT 0.0748125 0.36225 0.093122 0.38325 ;
  RECT 0.093122 0.18375 0.161437 0.202125 ;
  RECT 0.093122 0.36225 0.161437 0.38325 ;
  RECT 0.161437 0.18375 0.162094 0.202125 ;
  RECT 0.161437 0.202125 0.162094 0.2835 ;
  RECT 0.161437 0.36225 0.162094 0.38325 ;
  RECT 0.162094 0.18375 0.179812 0.202125 ;
  RECT 0.162094 0.202125 0.179812 0.2835 ;
  END
END XOR2_X1

END LIBRARY
#
# End of file
#
