# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2014, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *       NGLibraryCreator, Development_version_64 - build 201405271900        *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on us19.nangate.us for user Lucio Rech (lre).
# Local time is now Wed, 28 May 2014, 12:08:01.
# Main process id is 29163.

######Scaled from ocl15 by ChenlinShi 2022/1/6

VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.001 ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
  LAYER LEF58_PITCH STRING ;
  LAYER LEF58_GAP STRING ;
  LAYER LEF58_EOLKEEPOUT STRING ;
  LAYER LEF58_SPACING STRING ;
  LAYER LEF58_CORNERSPACING STRING ;
  LAYER LEF58_WIDTHTABLE STRING ;
  LAYER LEF58_CUTCLASS STRING ;
  LAYER LEF58_SPACINGTABLE STRING ;
  LAYER LEF58_ENCLOSURE STRING ;
  LAYER LEF58_RIGHTWAYONGRIDONLY STRING ;
  LAYER LEF58_RECTONLY STRING ;
END PROPERTYDEFINITIONS

LAYER nwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE PWELL ;" ;
END pwell



LAYER POLY
  TYPE MASTERSLICE ;
END POLY

LAYER ACT
  TYPE MASTERSLICE ;
END ACT

LAYER V0
  TYPE CUT ;
SPACING 0.010 ; 
WIDTH 0.022 ; 
END V0

LAYER M1
  TYPE ROUTING ;
SPACING 0.010 ; 
WIDTH 0.022 ; 
PITCH 0.032 0.032   ; 
  DIRECTION VERTICAL ;
OFFSET 0.000 0.016   ; 
END M1

LAYER V1
  TYPE CUT ;
SPACING 0.010 ; 
WIDTH 0.022 ; 

END V1

LAYER MINT1
  TYPE ROUTING ;
SPACING 0.018 ; 
WIDTH 0.024 ; 
PITCH 0.042 0.042   ; 
  DIRECTION HORIZONTAL ;
OFFSET 0.000 0.021   ; 
END MINT1

LAYER VINT1
  TYPE CUT ;
SPACING 0.016 ; 
WIDTH 0.016 ; 

END VINT1

LAYER MINT2
  TYPE ROUTING ;
SPACING 0.016 ; 
WIDTH 0.016 ; 
PITCH 0.032 0.032   ; 
  DIRECTION VERTICAL ;
OFFSET 0.000 0.016   ; 
END MINT2

LAYER VINT2
  TYPE CUT ;
SPACING 0.016 ; 
WIDTH 0.016 ; 

END VINT2

LAYER MINT3
  TYPE ROUTING ;
SPACING 0.016 ; 
WIDTH 0.016 ; 
PITCH 0.032 0.032   ; 
  DIRECTION HORIZONTAL ;
OFFSET 0.000 0.016   ; 
END MINT3

LAYER VINT3
  TYPE CUT ;
SPACING 0.024 ; 
WIDTH 0.016 ; 
END VINT3

LAYER MINT4
  TYPE ROUTING ;
SPACING 0.024 ; 
WIDTH 0.024 ; 
PITCH 0.048 0.048   ; 
  DIRECTION VERTICAL ;
OFFSET 0.000 0.024   ; 
END MINT4

LAYER VINT4
  TYPE CUT ;
SPACING 0.024 ; 
WIDTH 0.024 ; 

END VINT4

LAYER MINT5
  TYPE ROUTING ;
SPACING 0.024 ; 
WIDTH 0.024 ; 
PITCH 0.048 0.048   ; 
  DIRECTION HORIZONTAL ;
OFFSET 0.000 0.024   ; 
END MINT5

LAYER VINT5
  TYPE CUT ;
SPACING 0.040 ; 
WIDTH 0.024 ; 
END VINT5

LAYER MINT6
  TYPE ROUTING ;
SPACING 0.040 ; 
WIDTH 0.040 ; 
PITCH 0.080 0.080   ; 
  DIRECTION  VERTICAL ;
OFFSET 0.000 0.040   ; 
END MINT6

LAYER VINT6
  TYPE CUT ;
SPACING 0.040 ; 
WIDTH 0.040 ; 
END VINT6

LAYER MINT7
  TYPE ROUTING ;
SPACING 0.040 ; 
WIDTH 0.040 ; 
PITCH 0.080 0.080   ; 
  DIRECTION HORIZONTAL ;
OFFSET 0.000 0.040   ; 
END MINT7

LAYER VINT7
  TYPE CUT ;
SPACING 0.040 ; 
WIDTH 0.040 ; 
END VINT7

LAYER MINT8
  TYPE ROUTING ;
SPACING 0.040 ; 
WIDTH 0.040 ; 
PITCH 0.080 0.080   ; 
  DIRECTION VERTICAL ;
OFFSET 0.000 0.040   ; 
END MINT8


LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA V1_0 DEFAULT
  LAYER V1 ;
RECT -0.011 -0.011 0.011 0.011   ; 
  LAYER M1 ;
RECT -0.018 -0.018 0.018 0.018   ; 
  LAYER MINT1 ;
RECT -0.021 -0.021 0.021 0.021   ; 
END V1_0

VIA VINT1_0 DEFAULT
  LAYER VINT1 ;
RECT -0.008 -0.008 0.008 0.008   ; 
  LAYER MINT1 ;
RECT -0.021 -0.021 0.021 0.021   ; 
  LAYER MINT2 ;
RECT -0.014 -0.014 0.014 0.014   ; 
END VINT1_0

VIA VINT2_0 DEFAULT
  LAYER VINT2 ;
RECT -0.008 -0.008 0.008 0.008   ; 
  LAYER MINT2 ;
RECT -0.014 -0.014 0.014 0.014   ; 
  LAYER MINT3 ;
RECT -0.014 -0.014 0.014 0.014   ; 
END VINT2_0

VIA VINT3_0 DEFAULT
  LAYER VINT3 ;
RECT -0.008 -0.008 0.008 0.008   ; 
  LAYER MINT3 ;
RECT -0.014 -0.014 0.014 0.014   ; 
  LAYER MINT4 ;
RECT -0.021 -0.021 0.021 0.021   ; 
END VINT3_0

VIA VINT4_0 DEFAULT
  LAYER VINT4 ;
RECT -0.012 -0.012 0.012 0.012   ; 
  LAYER MINT4 ;
RECT -0.021 -0.021 0.021 0.021   ; 
  LAYER MINT5 ;
RECT -0.021 -0.021 0.021 0.021   ; 
END VINT4_0

VIA VINT5_0 DEFAULT
  LAYER VINT5 ;
RECT -0.012 -0.012 0.012 0.012   ; 
  LAYER MINT5 ;
RECT -0.021 -0.021 0.021 0.021   ; 
  LAYER MINT6 ;
RECT -0.034 -0.034 0.034 0.034   ; 
END VINT5_0

VIA VINT6_0 DEFAULT
  LAYER VINT6 ;
RECT -0.020 -0.020 0.020 0.020   ; 
  LAYER MINT6 ;
RECT -0.034 -0.034 0.034 0.034   ; 
  LAYER MINT7 ;
RECT -0.034 -0.034 0.034 0.034   ; 
END VINT6_0

VIA VINT7_0 DEFAULT
  LAYER VINT7 ;
RECT -0.020 -0.020 0.020 0.020   ; 
  LAYER MINT7 ;
RECT -0.034 -0.034 0.034 0.034   ; 
  LAYER MINT8 ;
RECT -0.034 -0.034 0.034 0.034   ; 
END VINT7_0

VIARULE Via1Array-0 GENERATE
  LAYER M1 ;
ENCLOSURE 0.024 0.000   ; 
  LAYER MINT1 ;
ENCLOSURE 0.027 0.000   ; 
  LAYER V1 ;
RECT -0.011 -0.011 0.011 0.011   ; 
SPACING 0.010 BY 0.010 ; 
END Via1Array-0

VIARULE Via1Array-1 GENERATE
  LAYER M1 ;
ENCLOSURE 0.000 0.024   ; 
  LAYER MINT1 ;
ENCLOSURE 0.000 0.027   ; 
  LAYER V1 ;
RECT -0.011 -0.011 0.011 0.011   ; 
SPACING 0.010 BY 0.010 ; 
END Via1Array-1

VIARULE Via1Array-2 GENERATE
  LAYER M1 ;
ENCLOSURE 0.024 0.000   ; 
  LAYER MINT1 ;
ENCLOSURE 0.000 0.027   ; 
  LAYER V1 ;
RECT -0.011 -0.011 0.011 0.011   ; 
SPACING 0.010 BY 0.010 ; 
END Via1Array-2

VIARULE Via1Array-3 GENERATE
  LAYER M1 ;
ENCLOSURE 0.000 0.024   ; 
  LAYER MINT1 ;
ENCLOSURE 0.027 0.000   ; 
  LAYER V1 ;
RECT -0.011 -0.011 0.011 0.011   ; 
SPACING 0.010 BY 0.010 ; 
END Via1Array-3

VIARULE Via1Array-4 GENERATE
  LAYER M1 ;
ENCLOSURE 0.021 0.002   ; 
  LAYER MINT1 ;
ENCLOSURE 0.024 0.002   ; 
  LAYER V1 ;
RECT -0.011 -0.011 0.011 0.011   ; 
SPACING 0.010 BY 0.010 ; 
END Via1Array-4

VIARULE Via1Array-5 GENERATE
  LAYER M1 ;
ENCLOSURE 0.002 0.021   ; 
  LAYER MINT1 ;
ENCLOSURE 0.002 0.024   ; 
  LAYER V1 ;
RECT -0.011 -0.011 0.011 0.011   ; 
SPACING 0.010 BY 0.010 ; 
END Via1Array-5

VIARULE Via1Array-6 GENERATE
  LAYER M1 ;
ENCLOSURE 0.002 0.021   ; 
  LAYER MINT1 ;
ENCLOSURE 0.024 0.002   ; 
  LAYER V1 ;
RECT -0.011 -0.011 0.011 0.011   ; 
SPACING 0.010 BY 0.010 ; 
END Via1Array-6

VIARULE Via1Array-7 GENERATE
  LAYER M1 ;
ENCLOSURE 0.021 0.002   ; 
  LAYER MINT1 ;
ENCLOSURE 0.002 0.024   ; 
  LAYER V1 ;
RECT -0.011 -0.011 0.011 0.011   ; 
SPACING 0.010 BY 0.010 ; 
END Via1Array-7

VIARULE Via2Array-0 GENERATE
  LAYER MINT2 ;
ENCLOSURE 0.018 0.000   ; 
  LAYER MINT3 ;
ENCLOSURE 0.018 0.000   ; 
  LAYER VINT2 ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.016 BY 0.016 ; 
END Via2Array-0

VIARULE Via2Array-1 GENERATE
  LAYER MINT2 ;
ENCLOSURE 0.000 0.018   ; 
  LAYER MINT3 ;
ENCLOSURE 0.000 0.018   ; 
  LAYER VINT2 ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.016 BY 0.016 ; 
END Via2Array-1

VIARULE Via2Array-2 GENERATE
  LAYER MINT2 ;
ENCLOSURE 0.018 0.000   ; 
  LAYER MINT3 ;
ENCLOSURE 0.000 0.018   ; 
  LAYER VINT2 ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.016 BY 0.016 ; 
END Via2Array-2

VIARULE Via2Array-3 GENERATE
  LAYER MINT2 ;
ENCLOSURE 0.000 0.018   ; 
  LAYER MINT3 ;
ENCLOSURE 0.018 0.000   ; 
  LAYER VINT2 ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.016 BY 0.016 ; 
END Via2Array-3

VIARULE Via2Array-4 GENERATE
  LAYER MINT2 ;
ENCLOSURE 0.016 0.001   ; 
  LAYER MINT3 ;
ENCLOSURE 0.016 0.001   ; 
  LAYER VINT2 ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.016 BY 0.016 ; 
END Via2Array-4

VIARULE Via2Array-5 GENERATE
  LAYER MINT2 ;
ENCLOSURE 0.001 0.016   ; 
  LAYER MINT3 ;
ENCLOSURE 0.001 0.016   ; 
  LAYER VINT2 ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.016 BY 0.016 ; 
END Via2Array-5

VIARULE Via2Array-6 GENERATE
  LAYER MINT2 ;
ENCLOSURE 0.001 0.016   ; 
  LAYER MINT3 ;
ENCLOSURE 0.016 0.001   ; 
  LAYER VINT2 ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.016 BY 0.016 ; 
END Via2Array-6

VIARULE Via2Array-7 GENERATE
  LAYER MINT2 ;
ENCLOSURE 0.016 0.001   ; 
  LAYER MINT3 ;
ENCLOSURE 0.001 0.016   ; 
  LAYER VINT2 ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.016 BY 0.016 ; 
END Via2Array-7

VIARULE Via3Array-0 GENERATE
  LAYER MINT3 ;
ENCLOSURE 0.018 0.000   ; 
  LAYER MINT4 ;
ENCLOSURE 0.027 0.000   ; 
  LAYER VINT3 ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.024 BY 0.024 ; 
END Via3Array-0

VIARULE Via3Array-1 GENERATE
  LAYER MINT3 ;
ENCLOSURE 0.000 0.018   ; 
  LAYER MINT4 ;
ENCLOSURE 0.000 0.027   ; 
  LAYER VINT3 ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.024 BY 0.024 ; 
END Via3Array-1

VIARULE Via3Array-2 GENERATE
  LAYER MINT3 ;
ENCLOSURE 0.018 0.000   ; 
  LAYER MINT4 ;
ENCLOSURE 0.000 0.027   ; 
  LAYER VINT3 ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.024 BY 0.024 ; 
END Via3Array-2

VIARULE Via3Array-3 GENERATE
  LAYER MINT3 ;
ENCLOSURE 0.000 0.018   ; 
  LAYER MINT4 ;
ENCLOSURE 0.027 0.000   ; 
  LAYER VINT3 ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.024 BY 0.024 ; 
END Via3Array-3

VIARULE Via3Array-4 GENERATE
  LAYER MINT3 ;
ENCLOSURE 0.016 0.001   ; 
  LAYER MINT4 ;
ENCLOSURE 0.024 0.002   ; 
  LAYER VINT3 ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.024 BY 0.024 ; 
END Via3Array-4

VIARULE Via3Array-5 GENERATE
  LAYER MINT3 ;
ENCLOSURE 0.001 0.016   ; 
  LAYER MINT4 ;
ENCLOSURE 0.002 0.024   ; 
  LAYER VINT3 ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.024 BY 0.024 ; 
END Via3Array-5

VIARULE Via3Array-6 GENERATE
  LAYER MINT3 ;
ENCLOSURE 0.001 0.016   ; 
  LAYER MINT4 ;
ENCLOSURE 0.024 0.002   ; 
  LAYER VINT3 ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.024 BY 0.024 ; 
END Via3Array-6

VIARULE Via3Array-7 GENERATE
  LAYER MINT3 ;
ENCLOSURE 0.016 0.001   ; 
  LAYER MINT4 ;
ENCLOSURE 0.002 0.024   ; 
  LAYER VINT3 ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.024 BY 0.024 ; 
END Via3Array-7

VIARULE Via4Array-0 GENERATE
  LAYER MINT4 ;
ENCLOSURE 0.027 0.000   ; 
  LAYER MINT5 ;
ENCLOSURE 0.027 0.000   ; 
  LAYER VINT4 ;
RECT -0.012 -0.012 0.012 0.012   ; 
SPACING 0.024 BY 0.024 ; 
END Via4Array-0

VIARULE Via4Array-1 GENERATE
  LAYER MINT4 ;
ENCLOSURE 0.000 0.027   ; 
  LAYER MINT5 ;
ENCLOSURE 0.000 0.027   ; 
  LAYER VINT4 ;
RECT -0.012 -0.012 0.012 0.012   ; 
SPACING 0.024 BY 0.024 ; 
END Via4Array-1

VIARULE Via4Array-2 GENERATE
  LAYER MINT4 ;
ENCLOSURE 0.027 0.000   ; 
  LAYER MINT5 ;
ENCLOSURE 0.000 0.027   ; 
  LAYER VINT4 ;
RECT -0.012 -0.012 0.012 0.012   ; 
SPACING 0.024 BY 0.024 ; 
END Via4Array-2

VIARULE Via4Array-3 GENERATE
  LAYER MINT4 ;
ENCLOSURE 0.000 0.027   ; 
  LAYER MINT5 ;
ENCLOSURE 0.027 0.000   ; 
  LAYER VINT4 ;
RECT -0.012 -0.012 0.012 0.012   ; 
SPACING 0.024 BY 0.024 ; 
END Via4Array-3

VIARULE Via4Array-4 GENERATE
  LAYER MINT4 ;
ENCLOSURE 0.024 0.002   ; 
  LAYER MINT5 ;
ENCLOSURE 0.024 0.002   ; 
  LAYER VINT4 ;
RECT -0.012 -0.012 0.012 0.012   ; 
SPACING 0.024 BY 0.024 ; 
END Via4Array-4

VIARULE Via4Array-5 GENERATE
  LAYER MINT4 ;
ENCLOSURE 0.002 0.024   ; 
  LAYER MINT5 ;
ENCLOSURE 0.002 0.024   ; 
  LAYER VINT4 ;
RECT -0.012 -0.012 0.012 0.012   ; 
SPACING 0.024 BY 0.024 ; 
END Via4Array-5

VIARULE Via4Array-6 GENERATE
  LAYER MINT4 ;
ENCLOSURE 0.002 0.024   ; 
  LAYER MINT5 ;
ENCLOSURE 0.024 0.002   ; 
  LAYER VINT4 ;
RECT -0.012 -0.012 0.012 0.012   ; 
SPACING 0.024 BY 0.024 ; 
END Via4Array-6

VIARULE Via4Array-7 GENERATE
  LAYER MINT4 ;
ENCLOSURE 0.024 0.002   ; 
  LAYER MINT5 ;
ENCLOSURE 0.002 0.024   ; 
  LAYER VINT4 ;
RECT -0.012 -0.012 0.012 0.012   ; 
SPACING 0.024 BY 0.024 ; 
END Via4Array-7

VIARULE Via5Array-0 GENERATE
  LAYER MINT5 ;
ENCLOSURE 0.027 0.000   ; 
  LAYER MINT6 ;
ENCLOSURE 0.046 0.000   ; 
  LAYER VINT5 ;
RECT -0.012 -0.012 0.012 0.012   ; 
SPACING 0.040 BY 0.040 ; 
END Via5Array-0

VIARULE Via5Array-1 GENERATE
  LAYER MINT5 ;
ENCLOSURE 0.000 0.027   ; 
  LAYER MINT6 ;
ENCLOSURE 0.000 0.046   ; 
  LAYER VINT5 ;
RECT -0.012 -0.012 0.012 0.012   ; 
SPACING 0.040 BY 0.040 ; 
END Via5Array-1

VIARULE Via5Array-2 GENERATE
  LAYER MINT5 ;
ENCLOSURE 0.027 0.000   ; 
  LAYER MINT6 ;
ENCLOSURE 0.000 0.046   ; 
  LAYER VINT5 ;
RECT -0.012 -0.012 0.012 0.012   ; 
SPACING 0.040 BY 0.040 ; 
END Via5Array-2

VIARULE Via5Array-3 GENERATE
  LAYER MINT5 ;
ENCLOSURE 0.000 0.027   ; 
  LAYER MINT6 ;
ENCLOSURE 0.046 0.000   ; 
  LAYER VINT5 ;
RECT -0.012 -0.012 0.012 0.012   ; 
SPACING 0.040 BY 0.040 ; 
END Via5Array-3

VIARULE Via5Array-4 GENERATE
  LAYER MINT5 ;
ENCLOSURE 0.024 0.002   ; 
  LAYER MINT6 ;
ENCLOSURE 0.040 0.003   ; 
  LAYER VINT5 ;
RECT -0.012 -0.012 0.012 0.012   ; 
SPACING 0.040 BY 0.040 ; 
END Via5Array-4

VIARULE Via5Array-5 GENERATE
  LAYER MINT5 ;
ENCLOSURE 0.002 0.024   ; 
  LAYER MINT6 ;
ENCLOSURE 0.003 0.040   ; 
  LAYER VINT5 ;
RECT -0.012 -0.012 0.012 0.012   ; 
SPACING 0.040 BY 0.040 ; 
END Via5Array-5

VIARULE Via5Array-6 GENERATE
  LAYER MINT5 ;
ENCLOSURE 0.002 0.024   ; 
  LAYER MINT6 ;
ENCLOSURE 0.040 0.003   ; 
  LAYER VINT5 ;
RECT -0.012 -0.012 0.012 0.012   ; 
SPACING 0.040 BY 0.040 ; 
END Via5Array-6

VIARULE Via5Array-7 GENERATE
  LAYER MINT5 ;
ENCLOSURE 0.024 0.002   ; 
  LAYER MINT6 ;
ENCLOSURE 0.003 0.040   ; 
  LAYER VINT5 ;
RECT -0.012 -0.012 0.012 0.012   ; 
SPACING 0.040 BY 0.040 ; 
END Via5Array-7

VIARULE Via6Array-0 GENERATE
  LAYER MINT6 ;
ENCLOSURE 0.046 0.000   ; 
  LAYER MINT7 ;
ENCLOSURE 0.046 0.000   ; 
  LAYER VINT6 ;
RECT -0.020 -0.020 0.020 0.020   ; 
SPACING 0.040 BY 0.040 ; 
END Via6Array-0

VIARULE Via6Array-1 GENERATE
  LAYER MINT6 ;
ENCLOSURE 0.000 0.004   ; 
  LAYER MINT7 ;
ENCLOSURE 0.000 0.004   ; 
  LAYER VINT6 ;
RECT -0.020 -0.020 0.020 0.020   ; 
SPACING 0.040 BY 0.040 ; 
END Via6Array-1

VIARULE Via6Array-2 GENERATE
  LAYER MINT6 ;
ENCLOSURE 0.046 0.000   ; 
  LAYER MINT7 ;
ENCLOSURE 0.000 0.046   ; 
  LAYER VINT6 ;
RECT -0.020 -0.020 0.020 0.020   ; 
SPACING 0.040 BY 0.040 ; 
END Via6Array-2

VIARULE Via6Array-3 GENERATE
  LAYER MINT6 ;
ENCLOSURE 0.000 0.046   ; 
  LAYER MINT7 ;
ENCLOSURE 0.046 0.000   ; 
  LAYER VINT6 ;
RECT -0.020 -0.020 0.020 0.020   ; 
SPACING 0.040 BY 0.040 ; 
END Via6Array-3

VIARULE Via6Array-4 GENERATE
  LAYER MINT6 ;
ENCLOSURE 0.040 0.003   ; 
  LAYER MINT7 ;
ENCLOSURE 0.040 0.003   ; 
  LAYER VINT6 ;
RECT -0.020 -0.020 0.020 0.020   ; 
SPACING 0.040 BY 0.040 ; 
END Via6Array-4

VIARULE Via6Array-5 GENERATE
  LAYER MINT6 ;
ENCLOSURE 0.003 0.040   ; 
  LAYER MINT7 ;
ENCLOSURE 0.003 0.040   ; 
  LAYER VINT6 ;
RECT -0.020 -0.020 0.020 0.020   ; 
SPACING 0.040 BY 0.040 ; 
END Via6Array-5

VIARULE Via6Array-6 GENERATE
  LAYER MINT6 ;
ENCLOSURE 0.003 0.040   ; 
  LAYER MINT7 ;
ENCLOSURE 0.040 0.003   ; 
  LAYER VINT6 ;
RECT -0.020 -0.020 0.020 0.020   ; 
SPACING 0.040 BY 0.040 ; 
END Via6Array-6

VIARULE Via6Array-7 GENERATE
  LAYER MINT6 ;
ENCLOSURE 0.040 0.003   ; 
  LAYER MINT7 ;
ENCLOSURE 0.003 0.040   ; 
  LAYER VINT6 ;
RECT -0.020 -0.020 0.020 0.020   ; 
SPACING 0.040 BY 0.040 ; 
END Via6Array-7

VIARULE Via7Array-0 GENERATE
  LAYER MINT7 ;
ENCLOSURE 0.046 0.000   ; 
  LAYER MINT8 ;
ENCLOSURE 0.046 0.000   ; 
  LAYER VINT7 ;
RECT -0.020 -0.020 0.020 0.020   ; 
SPACING 0.040 BY 0.040 ; 
END Via7Array-0

VIARULE Via7Array-1 GENERATE
  LAYER MINT7 ;
ENCLOSURE 0.000 0.004   ; 
  LAYER MINT8 ;
ENCLOSURE 0.000 0.004   ; 
  LAYER VINT7  ;
RECT -0.020 -0.020 0.020 0.020   ; 
SPACING 0.040 BY 0.040 ; 
END Via7Array-1

VIARULE Via7Array-2 GENERATE
  LAYER MINT7 ;
ENCLOSURE 0.046 0.000   ; 
  LAYER MINT8 ;
ENCLOSURE 0.000 0.046   ; 
  LAYER VINT7  ;
RECT -0.020 -0.020 0.020 0.020   ; 
SPACING 0.040 BY 0.040 ; 
END Via7Array-2

VIARULE Via7Array-3 GENERATE
  LAYER MINT7 ;
ENCLOSURE 0.000 0.046   ; 
  LAYER MINT8 ;
ENCLOSURE 0.046 0.000   ; 
  LAYER VINT7  ;
RECT -0.020 -0.020 0.020 0.020   ; 
SPACING 0.040 BY 0.040 ; 
END Via7Array-3

VIARULE Via7Array-4 GENERATE
  LAYER MINT7 ;
ENCLOSURE 0.040 0.003   ; 
  LAYER MINT8 ;
ENCLOSURE 0.040 0.003   ; 
  LAYER VINT7  ;
RECT -0.020 -0.020 0.020 0.020   ; 
SPACING 0.040 BY 0.040 ; 
END Via7Array-4

VIARULE Via7Array-5 GENERATE
  LAYER MINT7 ;
ENCLOSURE 0.003 0.040   ; 
  LAYER MINT8 ;
ENCLOSURE 0.003 0.040   ; 
  LAYER VINT7  ;
RECT -0.020 -0.020 0.020 0.020   ; 
SPACING 0.040 BY 0.040 ; 
END Via7Array-5

VIARULE Via7Array-6 GENERATE
  LAYER MINT7 ;
ENCLOSURE 0.003 0.040   ; 
  LAYER MINT8 ;
ENCLOSURE 0.040 0.003   ; 
  LAYER VINT7  ;
RECT -0.020 -0.020 0.020 0.020   ; 
SPACING 0.040 BY 0.040 ; 
END Via7Array-6

VIARULE Via7Array-7 GENERATE
  LAYER MINT7 ;
ENCLOSURE 0.040 0.003   ; 
  LAYER MINT8 ;
ENCLOSURE 0.003 0.040   ; 
  LAYER VINT7  ;
RECT -0.020 -0.020 0.020 0.020   ; 
SPACING 0.040 BY 0.040 ; 
END Via7Array-7

VIARULE Via8Array-0 GENERATE
  LAYER MINT1 ;
ENCLOSURE 0.027 0.000   ; 
  LAYER MINT2 ;
ENCLOSURE 0.018 0.000   ; 
  LAYER VINT1 ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.016 BY 0.016 ; 
END Via8Array-0

VIARULE Via8Array-1 GENERATE
  LAYER MINT1 ;
ENCLOSURE 0.000 0.027   ; 
  LAYER MINT2 ;
ENCLOSURE 0.000 0.018   ; 
  LAYER VINT1  ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.016 BY 0.016 ; 
END Via8Array-1

VIARULE Via8Array-2 GENERATE
  LAYER MINT1 ;
ENCLOSURE 0.027 0.000   ; 
  LAYER MINT2 ;
ENCLOSURE 0.000 0.018   ; 
  LAYER VINT1  ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.016 BY 0.016 ; 
END Via8Array-2

VIARULE Via8Array-3 GENERATE
  LAYER MINT1 ;
ENCLOSURE 0.000 0.027   ; 
  LAYER MINT2 ;
ENCLOSURE 0.018 0.000   ; 
  LAYER VINT1  ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.016 BY 0.016 ; 
END Via8Array-3

VIARULE Via8Array-4 GENERATE
  LAYER MINT1 ;
ENCLOSURE 0.024 0.002   ; 
  LAYER MINT2 ;
ENCLOSURE 0.016 0.001   ; 
  LAYER VINT1  ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.016 BY 0.016 ; 
END Via8Array-4

VIARULE Via8Array-5 GENERATE
  LAYER MINT1 ;
ENCLOSURE 0.002 0.024   ; 
  LAYER MINT2 ;
ENCLOSURE 0.001 0.016   ; 
  LAYER VINT1  ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.016 BY 0.016 ; 
END Via8Array-5

VIARULE Via8Array-6 GENERATE
  LAYER MINT1 ;
ENCLOSURE 0.002 0.024   ; 
  LAYER MINT2 ;
ENCLOSURE 0.016 0.001   ; 
  LAYER VINT1  ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.016 BY 0.016 ; 
END Via8Array-6

VIARULE Via8Array-7 GENERATE
  LAYER MINT1 ;
ENCLOSURE 0.024 0.002   ; 
  LAYER MINT2 ;
ENCLOSURE 0.001 0.016   ; 
  LAYER VINT1  ;
RECT -0.008 -0.008 0.008 0.008   ; 
SPACING 0.016 BY 0.016 ; 
END Via8Array-7

SPACING 
SAMENET M1 M1 0.010 ; 
SAMENET MINT2 MINT2 0.016 ; 
SAMENET MINT3 MINT3 0.016 ; 
SAMENET MINT4 MINT4 0.024 ; 
SAMENET MINT5 MINT5 0.024 ; 
SAMENET MINT6 MINT6 0.040 ; 
SAMENET MINT7 MINT7 0.040 ; 
SAMENET MINT8 MINT8 0.040 ; 
SAMENET V1 V1 0.010 ; 
SAMENET VINT2 VINT2 0.016 ; 
SAMENET VINT3 VINT3 0.024 ; 
SAMENET VINT4 VINT4 0.024 ; 
SAMENET VINT5 VINT5 0.040 ; 
SAMENET VINT6 VINT6 0.040 ; 
SAMENET VINT7 VINT7 0.040 ; 
SAMENET V1 VINT2 0.000 ; 
SAMENET VINT2 VINT3 0.000 ; 
SAMENET VINT3 VINT4 0.000 ; 
SAMENET VINT4 VINT5 0.000 ; 
SAMENET VINT5 VINT6 0.000 ; 
SAMENET VINT6 VINT7 0.000 ; 
END SPACING



END LIBRARY
#
# End of file
#
